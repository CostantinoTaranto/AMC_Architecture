
module AME_Architecture_expanded ( cMV0_in, cMV1_in, cMV2_in, START, CU_h, 
        CU_w, clk, RST, cREADY, VALID, eMV0_in, eMV1_in, eMV2_in, sixPar, 
        eIN_SEL, RefPel, CurPel, RADDR_RefCu_x, RADDR_RefCu_y, RADDR_CurCu_x, 
        RADDR_CurCu_y, MEM_RE, eREADY, eDONE, MV0_out, MV1_out, MV2_out, 
        cComp_EN, cDONE, eComp_EN, MVP0, MVP1, MVP2, CurSAD, D_Cur, 
        last_block_x, last_block_y, last_cand, Second_ready, CountTerm_OUT, 
        INTER_DATA_VALID_SET, INTER_DATA_VALID_RESET, ADD3_MVin_LE_fSET, 
        ADD3_MVin_LE_nSET, ADD3_MVin_LE_fRESET, LE_ab, SAD_tmp_RST, Comp_EN, 
        OUT_LE, CountTerm_EN, CandCount_CE, RF_in_RE, BestCand, MULT1_VALID, 
        ADD3_VALID, incrY, ADD3_MVin_LE, eCU_PS, eCU_NS );
  input [21:0] cMV0_in;
  input [21:0] cMV1_in;
  input [21:0] cMV2_in;
  input [6:0] CU_h;
  input [6:0] CU_w;
  input [21:0] eMV0_in;
  input [21:0] eMV1_in;
  input [21:0] eMV2_in;
  input [31:0] RefPel;
  input [31:0] CurPel;
  output [12:0] RADDR_RefCu_x;
  output [12:0] RADDR_RefCu_y;
  output [5:0] RADDR_CurCu_x;
  output [5:0] RADDR_CurCu_y;
  output [21:0] MV0_out;
  output [21:0] MV1_out;
  output [21:0] MV2_out;
  output [21:0] MVP0;
  output [21:0] MVP1;
  output [21:0] MVP2;
  output [17:0] CurSAD;
  output [27:0] D_Cur;
  output [4:0] eCU_PS;
  output [4:0] eCU_NS;
  input START, clk, RST, VALID, sixPar, eIN_SEL;
  output cREADY, MEM_RE, eREADY, eDONE, cComp_EN, cDONE, eComp_EN,
         last_block_x, last_block_y, last_cand, Second_ready, CountTerm_OUT,
         INTER_DATA_VALID_SET, INTER_DATA_VALID_RESET, ADD3_MVin_LE_fSET,
         ADD3_MVin_LE_nSET, ADD3_MVin_LE_fRESET, LE_ab, SAD_tmp_RST, Comp_EN,
         OUT_LE, CountTerm_EN, CandCount_CE, RF_in_RE, BestCand, MULT1_VALID,
         ADD3_VALID, incrY, ADD3_MVin_LE;
  wire   eComp_EN, ADD3_MVin_LE_nSET, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243,
         constructing_unit_CE_compEN_int, constructing_unit_cmd_SH_EN_int,
         constructing_unit_RST_int, constructing_unit_CNT_STOPcompEN_OUT_int,
         constructing_unit_CNT_compEN_OUT_int,
         constructing_unit_Control_Unit_n6, constructing_unit_Control_Unit_n4,
         constructing_unit_Control_Unit_n3, constructing_unit_Control_Unit_n2,
         constructing_unit_Control_Unit_n1, constructing_unit_Control_Unit_n16,
         constructing_unit_Control_Unit_n15,
         constructing_unit_Control_Unit_n14,
         constructing_unit_Control_Unit_n13,
         constructing_unit_Control_Unit_n12,
         constructing_unit_Control_Unit_n11,
         constructing_unit_Control_Unit_n10, constructing_unit_Control_Unit_n9,
         constructing_unit_Control_Unit_n8, constructing_unit_Control_Unit_n7,
         constructing_unit_Control_Unit_PS_0_,
         constructing_unit_Control_Unit_PS_1_,
         constructing_unit_Control_Unit_PS_2_,
         constructing_unit_Control_Unit_CNT_STOPcompEN_OUT_int,
         constructing_unit_Control_Unit_CNT_compEN_OUT_int,
         constructing_unit_Control_Unit_GOT_int,
         constructing_unit_Control_Unit_START_int,
         constructing_unit_Control_Unit_START_sampling_n1,
         constructing_unit_Control_Unit_GOT_sampling_n1,
         constructing_unit_Control_Unit_CNT_compEN_OUT_sampling_n1,
         constructing_unit_Control_Unit_CNT_STOPcompEN_OUT_sampling_n1,
         constructing_unit_Datapath_n76, constructing_unit_Datapath_n75,
         constructing_unit_Datapath_n74, constructing_unit_Datapath_n73,
         constructing_unit_Datapath_n72, constructing_unit_Datapath_n71,
         constructing_unit_Datapath_n70, constructing_unit_Datapath_n69,
         constructing_unit_Datapath_n68, constructing_unit_Datapath_n67,
         constructing_unit_Datapath_n66, constructing_unit_Datapath_n65,
         constructing_unit_Datapath_n64, constructing_unit_Datapath_n63,
         constructing_unit_Datapath_n62, constructing_unit_Datapath_n61,
         constructing_unit_Datapath_n60, constructing_unit_Datapath_n59,
         constructing_unit_Datapath_n58, constructing_unit_Datapath_n29,
         constructing_unit_Datapath_n28, constructing_unit_Datapath_n27,
         constructing_unit_Datapath_n26, constructing_unit_Datapath_n25,
         constructing_unit_Datapath_n24, constructing_unit_Datapath_n23,
         constructing_unit_Datapath_n22, constructing_unit_Datapath_n21,
         constructing_unit_Datapath_n20, constructing_unit_Datapath_n19,
         constructing_unit_Datapath_n18, constructing_unit_Datapath_n17,
         constructing_unit_Datapath_n16, constructing_unit_Datapath_n15,
         constructing_unit_Datapath_n14, constructing_unit_Datapath_n13,
         constructing_unit_Datapath_n12, constructing_unit_Datapath_n11,
         constructing_unit_Datapath_n10, constructing_unit_Datapath_n9,
         constructing_unit_Datapath_n8, constructing_unit_Datapath_n7,
         constructing_unit_Datapath_n6, constructing_unit_Datapath_n5,
         constructing_unit_Datapath_n4, constructing_unit_Datapath_n3,
         constructing_unit_Datapath_n2, constructing_unit_Datapath_n1,
         constructing_unit_Datapath_n57, constructing_unit_Datapath_n56,
         constructing_unit_Datapath_n55, constructing_unit_Datapath_n54,
         constructing_unit_Datapath_n53, constructing_unit_Datapath_n52,
         constructing_unit_Datapath_n51, constructing_unit_Datapath_n50,
         constructing_unit_Datapath_n49, constructing_unit_Datapath_n48,
         constructing_unit_Datapath_n47, constructing_unit_Datapath_n46,
         constructing_unit_Datapath_n45, constructing_unit_Datapath_n44,
         constructing_unit_Datapath_n43, constructing_unit_Datapath_n42,
         constructing_unit_Datapath_n41, constructing_unit_Datapath_n40,
         constructing_unit_Datapath_n39, constructing_unit_Datapath_n38,
         constructing_unit_Datapath_n37, constructing_unit_Datapath_n36,
         constructing_unit_Datapath_n35, constructing_unit_Datapath_n34,
         constructing_unit_Datapath_n33, constructing_unit_Datapath_n32,
         constructing_unit_Datapath_n31, constructing_unit_Datapath_n30,
         constructing_unit_Datapath_comp_out,
         constructing_unit_Datapath_comp_out_tmp,
         constructing_unit_Datapath_comp_out_d,
         constructing_unit_Datapath_D_D_0_, constructing_unit_Datapath_D_D_1_,
         constructing_unit_Datapath_D_D_2_, constructing_unit_Datapath_D_D_3_,
         constructing_unit_Datapath_D_D_4_, constructing_unit_Datapath_D_D_5_,
         constructing_unit_Datapath_D_D_6_, constructing_unit_Datapath_D_D_7_,
         constructing_unit_Datapath_D_D_8_, constructing_unit_Datapath_D_D_9_,
         constructing_unit_Datapath_D_D_10_,
         constructing_unit_Datapath_D_D_11_,
         constructing_unit_Datapath_D_D_12_,
         constructing_unit_Datapath_D_D_13_,
         constructing_unit_Datapath_D_D_14_,
         constructing_unit_Datapath_D_D_15_,
         constructing_unit_Datapath_D_D_16_,
         constructing_unit_Datapath_D_D_17_,
         constructing_unit_Datapath_D_D_18_,
         constructing_unit_Datapath_D_D_19_,
         constructing_unit_Datapath_D_D_20_,
         constructing_unit_Datapath_D_D_21_,
         constructing_unit_Datapath_D_D_22_,
         constructing_unit_Datapath_D_D_23_,
         constructing_unit_Datapath_D_D_24_,
         constructing_unit_Datapath_D_D_25_,
         constructing_unit_Datapath_D_D_26_,
         constructing_unit_Datapath_D_D_27_,
         constructing_unit_Datapath_UA_flag_int_0_,
         constructing_unit_Datapath_UA_flag_int_1_,
         constructing_unit_Datapath_UA_flag_int_2_,
         constructing_unit_Datapath_UA_flag_int_3_,
         constructing_unit_Datapath_UA_flag_int_4_,
         constructing_unit_Datapath_UA_flag_int_5_,
         constructing_unit_Datapath_UA_flag_int_6_,
         constructing_unit_Datapath_UA_flag_int_7_,
         constructing_unit_Datapath_UA_flag_int_8_,
         constructing_unit_Datapath_UA_flag_int_9_,
         constructing_unit_Datapath_UA_flag_int_10_,
         constructing_unit_Datapath_D_v_0_, constructing_unit_Datapath_D_v_1_,
         constructing_unit_Datapath_D_v_2_, constructing_unit_Datapath_D_v_3_,
         constructing_unit_Datapath_D_v_4_, constructing_unit_Datapath_D_v_5_,
         constructing_unit_Datapath_D_v_6_, constructing_unit_Datapath_D_v_7_,
         constructing_unit_Datapath_D_v_8_, constructing_unit_Datapath_D_v_9_,
         constructing_unit_Datapath_D_v_10_,
         constructing_unit_Datapath_D_v_11_,
         constructing_unit_Datapath_D_v_12_,
         constructing_unit_Datapath_D_v_13_,
         constructing_unit_Datapath_D_v_14_,
         constructing_unit_Datapath_MV2_int_v_1__0_,
         constructing_unit_Datapath_MV2_int_v_1__1_,
         constructing_unit_Datapath_MV2_int_v_1__2_,
         constructing_unit_Datapath_MV2_int_v_1__3_,
         constructing_unit_Datapath_MV2_int_v_1__4_,
         constructing_unit_Datapath_MV2_int_v_1__5_,
         constructing_unit_Datapath_MV2_int_v_1__6_,
         constructing_unit_Datapath_MV2_int_v_1__7_,
         constructing_unit_Datapath_MV2_int_v_1__8_,
         constructing_unit_Datapath_MV2_int_v_1__9_,
         constructing_unit_Datapath_MV2_int_v_1__10_,
         constructing_unit_Datapath_MV2_int_v_2__0_,
         constructing_unit_Datapath_MV2_int_v_2__1_,
         constructing_unit_Datapath_MV2_int_v_2__2_,
         constructing_unit_Datapath_MV2_int_v_2__3_,
         constructing_unit_Datapath_MV2_int_v_2__4_,
         constructing_unit_Datapath_MV2_int_v_2__5_,
         constructing_unit_Datapath_MV2_int_v_2__6_,
         constructing_unit_Datapath_MV2_int_v_2__7_,
         constructing_unit_Datapath_MV2_int_v_2__8_,
         constructing_unit_Datapath_MV2_int_v_2__9_,
         constructing_unit_Datapath_MV2_int_v_2__10_,
         constructing_unit_Datapath_MV2_int_v_3__0_,
         constructing_unit_Datapath_MV2_int_v_3__1_,
         constructing_unit_Datapath_MV2_int_v_3__2_,
         constructing_unit_Datapath_MV2_int_v_3__3_,
         constructing_unit_Datapath_MV2_int_v_3__4_,
         constructing_unit_Datapath_MV2_int_v_3__5_,
         constructing_unit_Datapath_MV2_int_v_3__6_,
         constructing_unit_Datapath_MV2_int_v_3__7_,
         constructing_unit_Datapath_MV2_int_v_3__8_,
         constructing_unit_Datapath_MV2_int_v_3__9_,
         constructing_unit_Datapath_MV2_int_v_3__10_,
         constructing_unit_Datapath_MV2_int_v_4__0_,
         constructing_unit_Datapath_MV2_int_v_4__1_,
         constructing_unit_Datapath_MV2_int_v_4__2_,
         constructing_unit_Datapath_MV2_int_v_4__3_,
         constructing_unit_Datapath_MV2_int_v_4__4_,
         constructing_unit_Datapath_MV2_int_v_4__5_,
         constructing_unit_Datapath_MV2_int_v_4__6_,
         constructing_unit_Datapath_MV2_int_v_4__7_,
         constructing_unit_Datapath_MV2_int_v_4__8_,
         constructing_unit_Datapath_MV2_int_v_4__9_,
         constructing_unit_Datapath_MV2_int_v_4__10_,
         constructing_unit_Datapath_MV2_int_v_5__0_,
         constructing_unit_Datapath_MV2_int_v_5__1_,
         constructing_unit_Datapath_MV2_int_v_5__2_,
         constructing_unit_Datapath_MV2_int_v_5__3_,
         constructing_unit_Datapath_MV2_int_v_5__4_,
         constructing_unit_Datapath_MV2_int_v_5__5_,
         constructing_unit_Datapath_MV2_int_v_5__6_,
         constructing_unit_Datapath_MV2_int_v_5__7_,
         constructing_unit_Datapath_MV2_int_v_5__8_,
         constructing_unit_Datapath_MV2_int_v_5__9_,
         constructing_unit_Datapath_MV2_int_v_5__10_,
         constructing_unit_Datapath_MV2_int_v_6__0_,
         constructing_unit_Datapath_MV2_int_v_6__1_,
         constructing_unit_Datapath_MV2_int_v_6__2_,
         constructing_unit_Datapath_MV2_int_v_6__3_,
         constructing_unit_Datapath_MV2_int_v_6__4_,
         constructing_unit_Datapath_MV2_int_v_6__5_,
         constructing_unit_Datapath_MV2_int_v_6__6_,
         constructing_unit_Datapath_MV2_int_v_6__7_,
         constructing_unit_Datapath_MV2_int_v_6__8_,
         constructing_unit_Datapath_MV2_int_v_6__9_,
         constructing_unit_Datapath_MV2_int_v_6__10_,
         constructing_unit_Datapath_MV2_int_v_7__0_,
         constructing_unit_Datapath_MV2_int_v_7__1_,
         constructing_unit_Datapath_MV2_int_v_7__2_,
         constructing_unit_Datapath_MV2_int_v_7__3_,
         constructing_unit_Datapath_MV2_int_v_7__4_,
         constructing_unit_Datapath_MV2_int_v_7__5_,
         constructing_unit_Datapath_MV2_int_v_7__6_,
         constructing_unit_Datapath_MV2_int_v_7__7_,
         constructing_unit_Datapath_MV2_int_v_7__8_,
         constructing_unit_Datapath_MV2_int_v_7__9_,
         constructing_unit_Datapath_MV2_int_v_7__10_,
         constructing_unit_Datapath_MV2_int_v_9__0_,
         constructing_unit_Datapath_MV2_int_v_9__1_,
         constructing_unit_Datapath_MV2_int_v_9__2_,
         constructing_unit_Datapath_MV2_int_v_9__3_,
         constructing_unit_Datapath_MV2_int_v_9__4_,
         constructing_unit_Datapath_MV2_int_v_9__5_,
         constructing_unit_Datapath_MV2_int_v_9__6_,
         constructing_unit_Datapath_MV2_int_v_9__7_,
         constructing_unit_Datapath_MV2_int_v_9__8_,
         constructing_unit_Datapath_MV2_int_v_9__9_,
         constructing_unit_Datapath_MV2_int_v_9__10_,
         constructing_unit_Datapath_MV2_int_v_10__0_,
         constructing_unit_Datapath_MV2_int_v_10__1_,
         constructing_unit_Datapath_MV2_int_v_10__2_,
         constructing_unit_Datapath_MV2_int_v_10__3_,
         constructing_unit_Datapath_MV2_int_v_10__4_,
         constructing_unit_Datapath_MV2_int_v_10__5_,
         constructing_unit_Datapath_MV2_int_v_10__6_,
         constructing_unit_Datapath_MV2_int_v_10__7_,
         constructing_unit_Datapath_MV2_int_v_10__8_,
         constructing_unit_Datapath_MV2_int_v_10__9_,
         constructing_unit_Datapath_MV2_int_v_10__10_,
         constructing_unit_Datapath_MV2_int_v_11__0_,
         constructing_unit_Datapath_MV2_int_v_11__1_,
         constructing_unit_Datapath_MV2_int_v_11__2_,
         constructing_unit_Datapath_MV2_int_v_11__3_,
         constructing_unit_Datapath_MV2_int_v_11__4_,
         constructing_unit_Datapath_MV2_int_v_11__5_,
         constructing_unit_Datapath_MV2_int_v_11__6_,
         constructing_unit_Datapath_MV2_int_v_11__7_,
         constructing_unit_Datapath_MV2_int_v_11__8_,
         constructing_unit_Datapath_MV2_int_v_11__9_,
         constructing_unit_Datapath_MV2_int_v_11__10_,
         constructing_unit_Datapath_MV2_int_v_12__0_,
         constructing_unit_Datapath_MV2_int_v_12__1_,
         constructing_unit_Datapath_MV2_int_v_12__2_,
         constructing_unit_Datapath_MV2_int_v_12__3_,
         constructing_unit_Datapath_MV2_int_v_12__4_,
         constructing_unit_Datapath_MV2_int_v_12__5_,
         constructing_unit_Datapath_MV2_int_v_12__6_,
         constructing_unit_Datapath_MV2_int_v_12__7_,
         constructing_unit_Datapath_MV2_int_v_12__8_,
         constructing_unit_Datapath_MV2_int_v_12__9_,
         constructing_unit_Datapath_MV2_int_v_12__10_,
         constructing_unit_Datapath_MV2_int_v_13__0_,
         constructing_unit_Datapath_MV2_int_v_13__1_,
         constructing_unit_Datapath_MV2_int_v_13__2_,
         constructing_unit_Datapath_MV2_int_v_13__3_,
         constructing_unit_Datapath_MV2_int_v_13__4_,
         constructing_unit_Datapath_MV2_int_v_13__5_,
         constructing_unit_Datapath_MV2_int_v_13__6_,
         constructing_unit_Datapath_MV2_int_v_13__7_,
         constructing_unit_Datapath_MV2_int_v_13__8_,
         constructing_unit_Datapath_MV2_int_v_13__9_,
         constructing_unit_Datapath_MV2_int_v_13__10_,
         constructing_unit_Datapath_MV1_int_h_1__0_,
         constructing_unit_Datapath_MV1_int_h_1__1_,
         constructing_unit_Datapath_MV1_int_h_1__2_,
         constructing_unit_Datapath_MV1_int_h_1__3_,
         constructing_unit_Datapath_MV1_int_h_1__4_,
         constructing_unit_Datapath_MV1_int_h_1__5_,
         constructing_unit_Datapath_MV1_int_h_1__6_,
         constructing_unit_Datapath_MV1_int_h_1__7_,
         constructing_unit_Datapath_MV1_int_h_1__8_,
         constructing_unit_Datapath_MV1_int_h_1__9_,
         constructing_unit_Datapath_MV1_int_h_1__10_,
         constructing_unit_Datapath_MV1_int_h_2__0_,
         constructing_unit_Datapath_MV1_int_h_2__1_,
         constructing_unit_Datapath_MV1_int_h_2__2_,
         constructing_unit_Datapath_MV1_int_h_2__3_,
         constructing_unit_Datapath_MV1_int_h_2__4_,
         constructing_unit_Datapath_MV1_int_h_2__5_,
         constructing_unit_Datapath_MV1_int_h_2__6_,
         constructing_unit_Datapath_MV1_int_h_2__7_,
         constructing_unit_Datapath_MV1_int_h_2__8_,
         constructing_unit_Datapath_MV1_int_h_2__9_,
         constructing_unit_Datapath_MV1_int_h_2__10_,
         constructing_unit_Datapath_MV1_int_h_3__0_,
         constructing_unit_Datapath_MV1_int_h_3__1_,
         constructing_unit_Datapath_MV1_int_h_3__2_,
         constructing_unit_Datapath_MV1_int_h_3__3_,
         constructing_unit_Datapath_MV1_int_h_3__4_,
         constructing_unit_Datapath_MV1_int_h_3__5_,
         constructing_unit_Datapath_MV1_int_h_3__6_,
         constructing_unit_Datapath_MV1_int_h_3__7_,
         constructing_unit_Datapath_MV1_int_h_3__8_,
         constructing_unit_Datapath_MV1_int_h_3__9_,
         constructing_unit_Datapath_MV1_int_h_3__10_,
         constructing_unit_Datapath_MV1_int_h_4__0_,
         constructing_unit_Datapath_MV1_int_h_4__1_,
         constructing_unit_Datapath_MV1_int_h_4__2_,
         constructing_unit_Datapath_MV1_int_h_4__3_,
         constructing_unit_Datapath_MV1_int_h_4__4_,
         constructing_unit_Datapath_MV1_int_h_4__5_,
         constructing_unit_Datapath_MV1_int_h_4__6_,
         constructing_unit_Datapath_MV1_int_h_4__7_,
         constructing_unit_Datapath_MV1_int_h_4__8_,
         constructing_unit_Datapath_MV1_int_h_4__9_,
         constructing_unit_Datapath_MV1_int_h_4__10_,
         constructing_unit_Datapath_MV1_int_h_5__0_,
         constructing_unit_Datapath_MV1_int_h_5__1_,
         constructing_unit_Datapath_MV1_int_h_5__2_,
         constructing_unit_Datapath_MV1_int_h_5__3_,
         constructing_unit_Datapath_MV1_int_h_5__4_,
         constructing_unit_Datapath_MV1_int_h_5__5_,
         constructing_unit_Datapath_MV1_int_h_5__6_,
         constructing_unit_Datapath_MV1_int_h_5__7_,
         constructing_unit_Datapath_MV1_int_h_5__8_,
         constructing_unit_Datapath_MV1_int_h_5__9_,
         constructing_unit_Datapath_MV1_int_h_5__10_,
         constructing_unit_Datapath_MV1_int_h_6__0_,
         constructing_unit_Datapath_MV1_int_h_6__1_,
         constructing_unit_Datapath_MV1_int_h_6__2_,
         constructing_unit_Datapath_MV1_int_h_6__3_,
         constructing_unit_Datapath_MV1_int_h_6__4_,
         constructing_unit_Datapath_MV1_int_h_6__5_,
         constructing_unit_Datapath_MV1_int_h_6__6_,
         constructing_unit_Datapath_MV1_int_h_6__7_,
         constructing_unit_Datapath_MV1_int_h_6__8_,
         constructing_unit_Datapath_MV1_int_h_6__9_,
         constructing_unit_Datapath_MV1_int_h_6__10_,
         constructing_unit_Datapath_MV1_int_h_7__0_,
         constructing_unit_Datapath_MV1_int_h_7__1_,
         constructing_unit_Datapath_MV1_int_h_7__2_,
         constructing_unit_Datapath_MV1_int_h_7__3_,
         constructing_unit_Datapath_MV1_int_h_7__4_,
         constructing_unit_Datapath_MV1_int_h_7__5_,
         constructing_unit_Datapath_MV1_int_h_7__6_,
         constructing_unit_Datapath_MV1_int_h_7__7_,
         constructing_unit_Datapath_MV1_int_h_7__8_,
         constructing_unit_Datapath_MV1_int_h_7__9_,
         constructing_unit_Datapath_MV1_int_h_7__10_,
         constructing_unit_Datapath_MV1_int_h_8__0_,
         constructing_unit_Datapath_MV1_int_h_8__1_,
         constructing_unit_Datapath_MV1_int_h_8__2_,
         constructing_unit_Datapath_MV1_int_h_8__3_,
         constructing_unit_Datapath_MV1_int_h_8__4_,
         constructing_unit_Datapath_MV1_int_h_8__5_,
         constructing_unit_Datapath_MV1_int_h_8__6_,
         constructing_unit_Datapath_MV1_int_h_8__7_,
         constructing_unit_Datapath_MV1_int_h_8__8_,
         constructing_unit_Datapath_MV1_int_h_8__9_,
         constructing_unit_Datapath_MV1_int_h_8__10_,
         constructing_unit_Datapath_MV1_int_h_9__0_,
         constructing_unit_Datapath_MV1_int_h_9__1_,
         constructing_unit_Datapath_MV1_int_h_9__2_,
         constructing_unit_Datapath_MV1_int_h_9__3_,
         constructing_unit_Datapath_MV1_int_h_9__4_,
         constructing_unit_Datapath_MV1_int_h_9__5_,
         constructing_unit_Datapath_MV1_int_h_9__6_,
         constructing_unit_Datapath_MV1_int_h_9__7_,
         constructing_unit_Datapath_MV1_int_h_9__8_,
         constructing_unit_Datapath_MV1_int_h_9__9_,
         constructing_unit_Datapath_MV1_int_h_9__10_,
         constructing_unit_Datapath_MV1_int_h_10__0_,
         constructing_unit_Datapath_MV1_int_h_10__1_,
         constructing_unit_Datapath_MV1_int_h_10__2_,
         constructing_unit_Datapath_MV1_int_h_10__3_,
         constructing_unit_Datapath_MV1_int_h_10__4_,
         constructing_unit_Datapath_MV1_int_h_10__5_,
         constructing_unit_Datapath_MV1_int_h_10__6_,
         constructing_unit_Datapath_MV1_int_h_10__7_,
         constructing_unit_Datapath_MV1_int_h_10__8_,
         constructing_unit_Datapath_MV1_int_h_10__9_,
         constructing_unit_Datapath_MV1_int_h_10__10_,
         constructing_unit_Datapath_MV1_int_h_11__0_,
         constructing_unit_Datapath_MV1_int_h_11__1_,
         constructing_unit_Datapath_MV1_int_h_11__2_,
         constructing_unit_Datapath_MV1_int_h_11__3_,
         constructing_unit_Datapath_MV1_int_h_11__4_,
         constructing_unit_Datapath_MV1_int_h_11__5_,
         constructing_unit_Datapath_MV1_int_h_11__6_,
         constructing_unit_Datapath_MV1_int_h_11__7_,
         constructing_unit_Datapath_MV1_int_h_11__8_,
         constructing_unit_Datapath_MV1_int_h_11__9_,
         constructing_unit_Datapath_MV1_int_h_11__10_,
         constructing_unit_Datapath_MV1_int_h_12__0_,
         constructing_unit_Datapath_MV1_int_h_12__1_,
         constructing_unit_Datapath_MV1_int_h_12__2_,
         constructing_unit_Datapath_MV1_int_h_12__3_,
         constructing_unit_Datapath_MV1_int_h_12__4_,
         constructing_unit_Datapath_MV1_int_h_12__5_,
         constructing_unit_Datapath_MV1_int_h_12__6_,
         constructing_unit_Datapath_MV1_int_h_12__7_,
         constructing_unit_Datapath_MV1_int_h_12__8_,
         constructing_unit_Datapath_MV1_int_h_12__9_,
         constructing_unit_Datapath_MV1_int_h_12__10_,
         constructing_unit_Datapath_MV1_int_h_13__0_,
         constructing_unit_Datapath_MV1_int_h_13__1_,
         constructing_unit_Datapath_MV1_int_h_13__2_,
         constructing_unit_Datapath_MV1_int_h_13__3_,
         constructing_unit_Datapath_MV1_int_h_13__4_,
         constructing_unit_Datapath_MV1_int_h_13__5_,
         constructing_unit_Datapath_MV1_int_h_13__6_,
         constructing_unit_Datapath_MV1_int_h_13__7_,
         constructing_unit_Datapath_MV1_int_h_13__8_,
         constructing_unit_Datapath_MV1_int_h_13__9_,
         constructing_unit_Datapath_MV1_int_h_13__10_,
         constructing_unit_Datapath_D_h_0_, constructing_unit_Datapath_D_h_1_,
         constructing_unit_Datapath_D_h_2_, constructing_unit_Datapath_D_h_3_,
         constructing_unit_Datapath_D_h_4_, constructing_unit_Datapath_D_h_5_,
         constructing_unit_Datapath_D_h_6_, constructing_unit_Datapath_D_h_7_,
         constructing_unit_Datapath_D_h_8_, constructing_unit_Datapath_D_h_9_,
         constructing_unit_Datapath_D_h_10_,
         constructing_unit_Datapath_D_h_11_,
         constructing_unit_Datapath_D_h_12_,
         constructing_unit_Datapath_D_h_13_,
         constructing_unit_Datapath_D_h_14_,
         constructing_unit_Datapath_MV2_int_h_1__0_,
         constructing_unit_Datapath_MV2_int_h_1__1_,
         constructing_unit_Datapath_MV2_int_h_1__2_,
         constructing_unit_Datapath_MV2_int_h_1__3_,
         constructing_unit_Datapath_MV2_int_h_1__4_,
         constructing_unit_Datapath_MV2_int_h_1__5_,
         constructing_unit_Datapath_MV2_int_h_1__6_,
         constructing_unit_Datapath_MV2_int_h_1__7_,
         constructing_unit_Datapath_MV2_int_h_1__8_,
         constructing_unit_Datapath_MV2_int_h_1__9_,
         constructing_unit_Datapath_MV2_int_h_1__10_,
         constructing_unit_Datapath_MV2_int_h_2__0_,
         constructing_unit_Datapath_MV2_int_h_2__1_,
         constructing_unit_Datapath_MV2_int_h_2__2_,
         constructing_unit_Datapath_MV2_int_h_2__3_,
         constructing_unit_Datapath_MV2_int_h_2__4_,
         constructing_unit_Datapath_MV2_int_h_2__5_,
         constructing_unit_Datapath_MV2_int_h_2__6_,
         constructing_unit_Datapath_MV2_int_h_2__7_,
         constructing_unit_Datapath_MV2_int_h_2__8_,
         constructing_unit_Datapath_MV2_int_h_2__9_,
         constructing_unit_Datapath_MV2_int_h_2__10_,
         constructing_unit_Datapath_MV2_int_h_3__0_,
         constructing_unit_Datapath_MV2_int_h_3__1_,
         constructing_unit_Datapath_MV2_int_h_3__2_,
         constructing_unit_Datapath_MV2_int_h_3__3_,
         constructing_unit_Datapath_MV2_int_h_3__4_,
         constructing_unit_Datapath_MV2_int_h_3__5_,
         constructing_unit_Datapath_MV2_int_h_3__6_,
         constructing_unit_Datapath_MV2_int_h_3__7_,
         constructing_unit_Datapath_MV2_int_h_3__8_,
         constructing_unit_Datapath_MV2_int_h_3__9_,
         constructing_unit_Datapath_MV2_int_h_3__10_,
         constructing_unit_Datapath_MV2_int_h_4__0_,
         constructing_unit_Datapath_MV2_int_h_4__1_,
         constructing_unit_Datapath_MV2_int_h_4__2_,
         constructing_unit_Datapath_MV2_int_h_4__3_,
         constructing_unit_Datapath_MV2_int_h_4__4_,
         constructing_unit_Datapath_MV2_int_h_4__5_,
         constructing_unit_Datapath_MV2_int_h_4__6_,
         constructing_unit_Datapath_MV2_int_h_4__7_,
         constructing_unit_Datapath_MV2_int_h_4__8_,
         constructing_unit_Datapath_MV2_int_h_4__9_,
         constructing_unit_Datapath_MV2_int_h_4__10_,
         constructing_unit_Datapath_MV2_int_h_5__0_,
         constructing_unit_Datapath_MV2_int_h_5__1_,
         constructing_unit_Datapath_MV2_int_h_5__2_,
         constructing_unit_Datapath_MV2_int_h_5__3_,
         constructing_unit_Datapath_MV2_int_h_5__4_,
         constructing_unit_Datapath_MV2_int_h_5__5_,
         constructing_unit_Datapath_MV2_int_h_5__6_,
         constructing_unit_Datapath_MV2_int_h_5__7_,
         constructing_unit_Datapath_MV2_int_h_5__8_,
         constructing_unit_Datapath_MV2_int_h_5__9_,
         constructing_unit_Datapath_MV2_int_h_5__10_,
         constructing_unit_Datapath_MV2_int_h_6__0_,
         constructing_unit_Datapath_MV2_int_h_6__1_,
         constructing_unit_Datapath_MV2_int_h_6__2_,
         constructing_unit_Datapath_MV2_int_h_6__3_,
         constructing_unit_Datapath_MV2_int_h_6__4_,
         constructing_unit_Datapath_MV2_int_h_6__5_,
         constructing_unit_Datapath_MV2_int_h_6__6_,
         constructing_unit_Datapath_MV2_int_h_6__7_,
         constructing_unit_Datapath_MV2_int_h_6__8_,
         constructing_unit_Datapath_MV2_int_h_6__9_,
         constructing_unit_Datapath_MV2_int_h_6__10_,
         constructing_unit_Datapath_MV2_int_h_7__0_,
         constructing_unit_Datapath_MV2_int_h_7__1_,
         constructing_unit_Datapath_MV2_int_h_7__2_,
         constructing_unit_Datapath_MV2_int_h_7__3_,
         constructing_unit_Datapath_MV2_int_h_7__4_,
         constructing_unit_Datapath_MV2_int_h_7__5_,
         constructing_unit_Datapath_MV2_int_h_7__6_,
         constructing_unit_Datapath_MV2_int_h_7__7_,
         constructing_unit_Datapath_MV2_int_h_7__8_,
         constructing_unit_Datapath_MV2_int_h_7__9_,
         constructing_unit_Datapath_MV2_int_h_7__10_,
         constructing_unit_Datapath_MV2_int_h_9__0_,
         constructing_unit_Datapath_MV2_int_h_9__1_,
         constructing_unit_Datapath_MV2_int_h_9__2_,
         constructing_unit_Datapath_MV2_int_h_9__3_,
         constructing_unit_Datapath_MV2_int_h_9__4_,
         constructing_unit_Datapath_MV2_int_h_9__5_,
         constructing_unit_Datapath_MV2_int_h_9__6_,
         constructing_unit_Datapath_MV2_int_h_9__7_,
         constructing_unit_Datapath_MV2_int_h_9__8_,
         constructing_unit_Datapath_MV2_int_h_9__9_,
         constructing_unit_Datapath_MV2_int_h_9__10_,
         constructing_unit_Datapath_MV2_int_h_10__0_,
         constructing_unit_Datapath_MV2_int_h_10__1_,
         constructing_unit_Datapath_MV2_int_h_10__2_,
         constructing_unit_Datapath_MV2_int_h_10__3_,
         constructing_unit_Datapath_MV2_int_h_10__4_,
         constructing_unit_Datapath_MV2_int_h_10__5_,
         constructing_unit_Datapath_MV2_int_h_10__6_,
         constructing_unit_Datapath_MV2_int_h_10__7_,
         constructing_unit_Datapath_MV2_int_h_10__8_,
         constructing_unit_Datapath_MV2_int_h_10__9_,
         constructing_unit_Datapath_MV2_int_h_10__10_,
         constructing_unit_Datapath_MV2_int_h_11__0_,
         constructing_unit_Datapath_MV2_int_h_11__1_,
         constructing_unit_Datapath_MV2_int_h_11__2_,
         constructing_unit_Datapath_MV2_int_h_11__3_,
         constructing_unit_Datapath_MV2_int_h_11__4_,
         constructing_unit_Datapath_MV2_int_h_11__5_,
         constructing_unit_Datapath_MV2_int_h_11__6_,
         constructing_unit_Datapath_MV2_int_h_11__7_,
         constructing_unit_Datapath_MV2_int_h_11__8_,
         constructing_unit_Datapath_MV2_int_h_11__9_,
         constructing_unit_Datapath_MV2_int_h_11__10_,
         constructing_unit_Datapath_MV2_int_h_12__0_,
         constructing_unit_Datapath_MV2_int_h_12__1_,
         constructing_unit_Datapath_MV2_int_h_12__2_,
         constructing_unit_Datapath_MV2_int_h_12__3_,
         constructing_unit_Datapath_MV2_int_h_12__4_,
         constructing_unit_Datapath_MV2_int_h_12__5_,
         constructing_unit_Datapath_MV2_int_h_12__6_,
         constructing_unit_Datapath_MV2_int_h_12__7_,
         constructing_unit_Datapath_MV2_int_h_12__8_,
         constructing_unit_Datapath_MV2_int_h_12__9_,
         constructing_unit_Datapath_MV2_int_h_12__10_,
         constructing_unit_Datapath_MV2_int_h_13__0_,
         constructing_unit_Datapath_MV2_int_h_13__1_,
         constructing_unit_Datapath_MV2_int_h_13__2_,
         constructing_unit_Datapath_MV2_int_h_13__3_,
         constructing_unit_Datapath_MV2_int_h_13__4_,
         constructing_unit_Datapath_MV2_int_h_13__5_,
         constructing_unit_Datapath_MV2_int_h_13__6_,
         constructing_unit_Datapath_MV2_int_h_13__7_,
         constructing_unit_Datapath_MV2_int_h_13__8_,
         constructing_unit_Datapath_MV2_int_h_13__9_,
         constructing_unit_Datapath_MV2_int_h_13__10_,
         constructing_unit_Datapath_MV0_int_h_1__0_,
         constructing_unit_Datapath_MV0_int_h_1__1_,
         constructing_unit_Datapath_MV0_int_h_1__2_,
         constructing_unit_Datapath_MV0_int_h_1__3_,
         constructing_unit_Datapath_MV0_int_h_1__4_,
         constructing_unit_Datapath_MV0_int_h_1__5_,
         constructing_unit_Datapath_MV0_int_h_1__6_,
         constructing_unit_Datapath_MV0_int_h_1__7_,
         constructing_unit_Datapath_MV0_int_h_1__8_,
         constructing_unit_Datapath_MV0_int_h_1__9_,
         constructing_unit_Datapath_MV0_int_h_1__10_,
         constructing_unit_Datapath_MV0_int_h_2__0_,
         constructing_unit_Datapath_MV0_int_h_2__1_,
         constructing_unit_Datapath_MV0_int_h_2__2_,
         constructing_unit_Datapath_MV0_int_h_2__3_,
         constructing_unit_Datapath_MV0_int_h_2__4_,
         constructing_unit_Datapath_MV0_int_h_2__5_,
         constructing_unit_Datapath_MV0_int_h_2__6_,
         constructing_unit_Datapath_MV0_int_h_2__7_,
         constructing_unit_Datapath_MV0_int_h_2__8_,
         constructing_unit_Datapath_MV0_int_h_2__9_,
         constructing_unit_Datapath_MV0_int_h_2__10_,
         constructing_unit_Datapath_MV0_int_h_3__0_,
         constructing_unit_Datapath_MV0_int_h_3__1_,
         constructing_unit_Datapath_MV0_int_h_3__2_,
         constructing_unit_Datapath_MV0_int_h_3__3_,
         constructing_unit_Datapath_MV0_int_h_3__4_,
         constructing_unit_Datapath_MV0_int_h_3__5_,
         constructing_unit_Datapath_MV0_int_h_3__6_,
         constructing_unit_Datapath_MV0_int_h_3__7_,
         constructing_unit_Datapath_MV0_int_h_3__8_,
         constructing_unit_Datapath_MV0_int_h_3__9_,
         constructing_unit_Datapath_MV0_int_h_3__10_,
         constructing_unit_Datapath_MV0_int_h_4__0_,
         constructing_unit_Datapath_MV0_int_h_4__1_,
         constructing_unit_Datapath_MV0_int_h_4__2_,
         constructing_unit_Datapath_MV0_int_h_4__3_,
         constructing_unit_Datapath_MV0_int_h_4__4_,
         constructing_unit_Datapath_MV0_int_h_4__5_,
         constructing_unit_Datapath_MV0_int_h_4__6_,
         constructing_unit_Datapath_MV0_int_h_4__7_,
         constructing_unit_Datapath_MV0_int_h_4__8_,
         constructing_unit_Datapath_MV0_int_h_4__9_,
         constructing_unit_Datapath_MV0_int_h_4__10_,
         constructing_unit_Datapath_MV0_int_h_5__0_,
         constructing_unit_Datapath_MV0_int_h_5__1_,
         constructing_unit_Datapath_MV0_int_h_5__2_,
         constructing_unit_Datapath_MV0_int_h_5__3_,
         constructing_unit_Datapath_MV0_int_h_5__4_,
         constructing_unit_Datapath_MV0_int_h_5__5_,
         constructing_unit_Datapath_MV0_int_h_5__6_,
         constructing_unit_Datapath_MV0_int_h_5__7_,
         constructing_unit_Datapath_MV0_int_h_5__8_,
         constructing_unit_Datapath_MV0_int_h_5__9_,
         constructing_unit_Datapath_MV0_int_h_5__10_,
         constructing_unit_Datapath_MV0_int_h_6__0_,
         constructing_unit_Datapath_MV0_int_h_6__1_,
         constructing_unit_Datapath_MV0_int_h_6__2_,
         constructing_unit_Datapath_MV0_int_h_6__3_,
         constructing_unit_Datapath_MV0_int_h_6__4_,
         constructing_unit_Datapath_MV0_int_h_6__5_,
         constructing_unit_Datapath_MV0_int_h_6__6_,
         constructing_unit_Datapath_MV0_int_h_6__7_,
         constructing_unit_Datapath_MV0_int_h_6__8_,
         constructing_unit_Datapath_MV0_int_h_6__9_,
         constructing_unit_Datapath_MV0_int_h_6__10_,
         constructing_unit_Datapath_MV0_int_h_8__0_,
         constructing_unit_Datapath_MV0_int_h_8__1_,
         constructing_unit_Datapath_MV0_int_h_8__2_,
         constructing_unit_Datapath_MV0_int_h_8__3_,
         constructing_unit_Datapath_MV0_int_h_8__4_,
         constructing_unit_Datapath_MV0_int_h_8__5_,
         constructing_unit_Datapath_MV0_int_h_8__6_,
         constructing_unit_Datapath_MV0_int_h_8__7_,
         constructing_unit_Datapath_MV0_int_h_8__8_,
         constructing_unit_Datapath_MV0_int_h_8__9_,
         constructing_unit_Datapath_MV0_int_h_8__10_,
         constructing_unit_Datapath_MV0_int_h_9__0_,
         constructing_unit_Datapath_MV0_int_h_9__1_,
         constructing_unit_Datapath_MV0_int_h_9__2_,
         constructing_unit_Datapath_MV0_int_h_9__3_,
         constructing_unit_Datapath_MV0_int_h_9__4_,
         constructing_unit_Datapath_MV0_int_h_9__5_,
         constructing_unit_Datapath_MV0_int_h_9__6_,
         constructing_unit_Datapath_MV0_int_h_9__7_,
         constructing_unit_Datapath_MV0_int_h_9__8_,
         constructing_unit_Datapath_MV0_int_h_9__9_,
         constructing_unit_Datapath_MV0_int_h_9__10_,
         constructing_unit_Datapath_MV0_int_h_10__0_,
         constructing_unit_Datapath_MV0_int_h_10__1_,
         constructing_unit_Datapath_MV0_int_h_10__2_,
         constructing_unit_Datapath_MV0_int_h_10__3_,
         constructing_unit_Datapath_MV0_int_h_10__4_,
         constructing_unit_Datapath_MV0_int_h_10__5_,
         constructing_unit_Datapath_MV0_int_h_10__6_,
         constructing_unit_Datapath_MV0_int_h_10__7_,
         constructing_unit_Datapath_MV0_int_h_10__8_,
         constructing_unit_Datapath_MV0_int_h_10__9_,
         constructing_unit_Datapath_MV0_int_h_10__10_,
         constructing_unit_Datapath_MV0_int_h_11__0_,
         constructing_unit_Datapath_MV0_int_h_11__1_,
         constructing_unit_Datapath_MV0_int_h_11__2_,
         constructing_unit_Datapath_MV0_int_h_11__3_,
         constructing_unit_Datapath_MV0_int_h_11__4_,
         constructing_unit_Datapath_MV0_int_h_11__5_,
         constructing_unit_Datapath_MV0_int_h_11__6_,
         constructing_unit_Datapath_MV0_int_h_11__7_,
         constructing_unit_Datapath_MV0_int_h_11__8_,
         constructing_unit_Datapath_MV0_int_h_11__9_,
         constructing_unit_Datapath_MV0_int_h_11__10_,
         constructing_unit_Datapath_MV0_int_h_12__0_,
         constructing_unit_Datapath_MV0_int_h_12__1_,
         constructing_unit_Datapath_MV0_int_h_12__2_,
         constructing_unit_Datapath_MV0_int_h_12__3_,
         constructing_unit_Datapath_MV0_int_h_12__4_,
         constructing_unit_Datapath_MV0_int_h_12__5_,
         constructing_unit_Datapath_MV0_int_h_12__6_,
         constructing_unit_Datapath_MV0_int_h_12__7_,
         constructing_unit_Datapath_MV0_int_h_12__8_,
         constructing_unit_Datapath_MV0_int_h_12__9_,
         constructing_unit_Datapath_MV0_int_h_12__10_,
         constructing_unit_Datapath_MV0_int_h_13__0_,
         constructing_unit_Datapath_MV0_int_h_13__1_,
         constructing_unit_Datapath_MV0_int_h_13__2_,
         constructing_unit_Datapath_MV0_int_h_13__3_,
         constructing_unit_Datapath_MV0_int_h_13__4_,
         constructing_unit_Datapath_MV0_int_h_13__5_,
         constructing_unit_Datapath_MV0_int_h_13__6_,
         constructing_unit_Datapath_MV0_int_h_13__7_,
         constructing_unit_Datapath_MV0_int_h_13__8_,
         constructing_unit_Datapath_MV0_int_h_13__9_,
         constructing_unit_Datapath_MV0_int_h_13__10_,
         constructing_unit_Datapath_SH_cmd_int_0_,
         constructing_unit_Datapath_SH_cmd_int_1_,
         constructing_unit_Datapath_SH_cmd_int_2_,
         constructing_unit_Datapath_MV0_int_v_1__0_,
         constructing_unit_Datapath_MV0_int_v_1__1_,
         constructing_unit_Datapath_MV0_int_v_1__2_,
         constructing_unit_Datapath_MV0_int_v_1__3_,
         constructing_unit_Datapath_MV0_int_v_1__4_,
         constructing_unit_Datapath_MV0_int_v_1__5_,
         constructing_unit_Datapath_MV0_int_v_1__6_,
         constructing_unit_Datapath_MV0_int_v_1__7_,
         constructing_unit_Datapath_MV0_int_v_1__8_,
         constructing_unit_Datapath_MV0_int_v_1__9_,
         constructing_unit_Datapath_MV0_int_v_1__10_,
         constructing_unit_Datapath_MV0_int_v_2__0_,
         constructing_unit_Datapath_MV0_int_v_2__1_,
         constructing_unit_Datapath_MV0_int_v_2__2_,
         constructing_unit_Datapath_MV0_int_v_2__3_,
         constructing_unit_Datapath_MV0_int_v_2__4_,
         constructing_unit_Datapath_MV0_int_v_2__5_,
         constructing_unit_Datapath_MV0_int_v_2__6_,
         constructing_unit_Datapath_MV0_int_v_2__7_,
         constructing_unit_Datapath_MV0_int_v_2__8_,
         constructing_unit_Datapath_MV0_int_v_2__9_,
         constructing_unit_Datapath_MV0_int_v_2__10_,
         constructing_unit_Datapath_MV0_int_v_3__0_,
         constructing_unit_Datapath_MV0_int_v_3__1_,
         constructing_unit_Datapath_MV0_int_v_3__2_,
         constructing_unit_Datapath_MV0_int_v_3__3_,
         constructing_unit_Datapath_MV0_int_v_3__4_,
         constructing_unit_Datapath_MV0_int_v_3__5_,
         constructing_unit_Datapath_MV0_int_v_3__6_,
         constructing_unit_Datapath_MV0_int_v_3__7_,
         constructing_unit_Datapath_MV0_int_v_3__8_,
         constructing_unit_Datapath_MV0_int_v_3__9_,
         constructing_unit_Datapath_MV0_int_v_3__10_,
         constructing_unit_Datapath_MV0_int_v_4__0_,
         constructing_unit_Datapath_MV0_int_v_4__1_,
         constructing_unit_Datapath_MV0_int_v_4__2_,
         constructing_unit_Datapath_MV0_int_v_4__3_,
         constructing_unit_Datapath_MV0_int_v_4__4_,
         constructing_unit_Datapath_MV0_int_v_4__5_,
         constructing_unit_Datapath_MV0_int_v_4__6_,
         constructing_unit_Datapath_MV0_int_v_4__7_,
         constructing_unit_Datapath_MV0_int_v_4__8_,
         constructing_unit_Datapath_MV0_int_v_4__9_,
         constructing_unit_Datapath_MV0_int_v_4__10_,
         constructing_unit_Datapath_MV0_int_v_5__0_,
         constructing_unit_Datapath_MV0_int_v_5__1_,
         constructing_unit_Datapath_MV0_int_v_5__2_,
         constructing_unit_Datapath_MV0_int_v_5__3_,
         constructing_unit_Datapath_MV0_int_v_5__4_,
         constructing_unit_Datapath_MV0_int_v_5__5_,
         constructing_unit_Datapath_MV0_int_v_5__6_,
         constructing_unit_Datapath_MV0_int_v_5__7_,
         constructing_unit_Datapath_MV0_int_v_5__8_,
         constructing_unit_Datapath_MV0_int_v_5__9_,
         constructing_unit_Datapath_MV0_int_v_5__10_,
         constructing_unit_Datapath_MV0_int_v_6__0_,
         constructing_unit_Datapath_MV0_int_v_6__1_,
         constructing_unit_Datapath_MV0_int_v_6__2_,
         constructing_unit_Datapath_MV0_int_v_6__3_,
         constructing_unit_Datapath_MV0_int_v_6__4_,
         constructing_unit_Datapath_MV0_int_v_6__5_,
         constructing_unit_Datapath_MV0_int_v_6__6_,
         constructing_unit_Datapath_MV0_int_v_6__7_,
         constructing_unit_Datapath_MV0_int_v_6__8_,
         constructing_unit_Datapath_MV0_int_v_6__9_,
         constructing_unit_Datapath_MV0_int_v_6__10_,
         constructing_unit_Datapath_MV0_int_v_8__0_,
         constructing_unit_Datapath_MV0_int_v_8__1_,
         constructing_unit_Datapath_MV0_int_v_8__2_,
         constructing_unit_Datapath_MV0_int_v_8__3_,
         constructing_unit_Datapath_MV0_int_v_8__4_,
         constructing_unit_Datapath_MV0_int_v_8__5_,
         constructing_unit_Datapath_MV0_int_v_8__6_,
         constructing_unit_Datapath_MV0_int_v_8__7_,
         constructing_unit_Datapath_MV0_int_v_8__8_,
         constructing_unit_Datapath_MV0_int_v_8__9_,
         constructing_unit_Datapath_MV0_int_v_8__10_,
         constructing_unit_Datapath_MV0_int_v_9__0_,
         constructing_unit_Datapath_MV0_int_v_9__1_,
         constructing_unit_Datapath_MV0_int_v_9__2_,
         constructing_unit_Datapath_MV0_int_v_9__3_,
         constructing_unit_Datapath_MV0_int_v_9__4_,
         constructing_unit_Datapath_MV0_int_v_9__5_,
         constructing_unit_Datapath_MV0_int_v_9__6_,
         constructing_unit_Datapath_MV0_int_v_9__7_,
         constructing_unit_Datapath_MV0_int_v_9__8_,
         constructing_unit_Datapath_MV0_int_v_9__9_,
         constructing_unit_Datapath_MV0_int_v_9__10_,
         constructing_unit_Datapath_MV0_int_v_10__0_,
         constructing_unit_Datapath_MV0_int_v_10__1_,
         constructing_unit_Datapath_MV0_int_v_10__2_,
         constructing_unit_Datapath_MV0_int_v_10__3_,
         constructing_unit_Datapath_MV0_int_v_10__4_,
         constructing_unit_Datapath_MV0_int_v_10__5_,
         constructing_unit_Datapath_MV0_int_v_10__6_,
         constructing_unit_Datapath_MV0_int_v_10__7_,
         constructing_unit_Datapath_MV0_int_v_10__8_,
         constructing_unit_Datapath_MV0_int_v_10__9_,
         constructing_unit_Datapath_MV0_int_v_10__10_,
         constructing_unit_Datapath_MV0_int_v_11__0_,
         constructing_unit_Datapath_MV0_int_v_11__1_,
         constructing_unit_Datapath_MV0_int_v_11__2_,
         constructing_unit_Datapath_MV0_int_v_11__3_,
         constructing_unit_Datapath_MV0_int_v_11__4_,
         constructing_unit_Datapath_MV0_int_v_11__5_,
         constructing_unit_Datapath_MV0_int_v_11__6_,
         constructing_unit_Datapath_MV0_int_v_11__7_,
         constructing_unit_Datapath_MV0_int_v_11__8_,
         constructing_unit_Datapath_MV0_int_v_11__9_,
         constructing_unit_Datapath_MV0_int_v_11__10_,
         constructing_unit_Datapath_MV0_int_v_12__0_,
         constructing_unit_Datapath_MV0_int_v_12__1_,
         constructing_unit_Datapath_MV0_int_v_12__2_,
         constructing_unit_Datapath_MV0_int_v_12__3_,
         constructing_unit_Datapath_MV0_int_v_12__4_,
         constructing_unit_Datapath_MV0_int_v_12__5_,
         constructing_unit_Datapath_MV0_int_v_12__6_,
         constructing_unit_Datapath_MV0_int_v_12__7_,
         constructing_unit_Datapath_MV0_int_v_12__8_,
         constructing_unit_Datapath_MV0_int_v_12__9_,
         constructing_unit_Datapath_MV0_int_v_12__10_,
         constructing_unit_Datapath_MV0_int_v_13__0_,
         constructing_unit_Datapath_MV0_int_v_13__1_,
         constructing_unit_Datapath_MV0_int_v_13__2_,
         constructing_unit_Datapath_MV0_int_v_13__3_,
         constructing_unit_Datapath_MV0_int_v_13__4_,
         constructing_unit_Datapath_MV0_int_v_13__5_,
         constructing_unit_Datapath_MV0_int_v_13__6_,
         constructing_unit_Datapath_MV0_int_v_13__7_,
         constructing_unit_Datapath_MV0_int_v_13__8_,
         constructing_unit_Datapath_MV0_int_v_13__9_,
         constructing_unit_Datapath_MV0_int_v_13__10_,
         constructing_unit_Datapath_MV1_int_v_1__0_,
         constructing_unit_Datapath_MV1_int_v_1__1_,
         constructing_unit_Datapath_MV1_int_v_1__2_,
         constructing_unit_Datapath_MV1_int_v_1__3_,
         constructing_unit_Datapath_MV1_int_v_1__4_,
         constructing_unit_Datapath_MV1_int_v_1__5_,
         constructing_unit_Datapath_MV1_int_v_1__6_,
         constructing_unit_Datapath_MV1_int_v_1__7_,
         constructing_unit_Datapath_MV1_int_v_1__8_,
         constructing_unit_Datapath_MV1_int_v_1__9_,
         constructing_unit_Datapath_MV1_int_v_1__10_,
         constructing_unit_Datapath_MV1_int_v_2__0_,
         constructing_unit_Datapath_MV1_int_v_2__1_,
         constructing_unit_Datapath_MV1_int_v_2__2_,
         constructing_unit_Datapath_MV1_int_v_2__3_,
         constructing_unit_Datapath_MV1_int_v_2__4_,
         constructing_unit_Datapath_MV1_int_v_2__5_,
         constructing_unit_Datapath_MV1_int_v_2__6_,
         constructing_unit_Datapath_MV1_int_v_2__7_,
         constructing_unit_Datapath_MV1_int_v_2__8_,
         constructing_unit_Datapath_MV1_int_v_2__9_,
         constructing_unit_Datapath_MV1_int_v_2__10_,
         constructing_unit_Datapath_MV1_int_v_3__0_,
         constructing_unit_Datapath_MV1_int_v_3__1_,
         constructing_unit_Datapath_MV1_int_v_3__2_,
         constructing_unit_Datapath_MV1_int_v_3__3_,
         constructing_unit_Datapath_MV1_int_v_3__4_,
         constructing_unit_Datapath_MV1_int_v_3__5_,
         constructing_unit_Datapath_MV1_int_v_3__6_,
         constructing_unit_Datapath_MV1_int_v_3__7_,
         constructing_unit_Datapath_MV1_int_v_3__8_,
         constructing_unit_Datapath_MV1_int_v_3__9_,
         constructing_unit_Datapath_MV1_int_v_3__10_,
         constructing_unit_Datapath_MV1_int_v_4__0_,
         constructing_unit_Datapath_MV1_int_v_4__1_,
         constructing_unit_Datapath_MV1_int_v_4__2_,
         constructing_unit_Datapath_MV1_int_v_4__3_,
         constructing_unit_Datapath_MV1_int_v_4__4_,
         constructing_unit_Datapath_MV1_int_v_4__5_,
         constructing_unit_Datapath_MV1_int_v_4__6_,
         constructing_unit_Datapath_MV1_int_v_4__7_,
         constructing_unit_Datapath_MV1_int_v_4__8_,
         constructing_unit_Datapath_MV1_int_v_4__9_,
         constructing_unit_Datapath_MV1_int_v_4__10_,
         constructing_unit_Datapath_MV1_int_v_5__0_,
         constructing_unit_Datapath_MV1_int_v_5__1_,
         constructing_unit_Datapath_MV1_int_v_5__2_,
         constructing_unit_Datapath_MV1_int_v_5__3_,
         constructing_unit_Datapath_MV1_int_v_5__4_,
         constructing_unit_Datapath_MV1_int_v_5__5_,
         constructing_unit_Datapath_MV1_int_v_5__6_,
         constructing_unit_Datapath_MV1_int_v_5__7_,
         constructing_unit_Datapath_MV1_int_v_5__8_,
         constructing_unit_Datapath_MV1_int_v_5__9_,
         constructing_unit_Datapath_MV1_int_v_5__10_,
         constructing_unit_Datapath_MV1_int_v_6__0_,
         constructing_unit_Datapath_MV1_int_v_6__1_,
         constructing_unit_Datapath_MV1_int_v_6__2_,
         constructing_unit_Datapath_MV1_int_v_6__3_,
         constructing_unit_Datapath_MV1_int_v_6__4_,
         constructing_unit_Datapath_MV1_int_v_6__5_,
         constructing_unit_Datapath_MV1_int_v_6__6_,
         constructing_unit_Datapath_MV1_int_v_6__7_,
         constructing_unit_Datapath_MV1_int_v_6__8_,
         constructing_unit_Datapath_MV1_int_v_6__9_,
         constructing_unit_Datapath_MV1_int_v_6__10_,
         constructing_unit_Datapath_MV1_int_v_7__0_,
         constructing_unit_Datapath_MV1_int_v_7__1_,
         constructing_unit_Datapath_MV1_int_v_7__2_,
         constructing_unit_Datapath_MV1_int_v_7__3_,
         constructing_unit_Datapath_MV1_int_v_7__4_,
         constructing_unit_Datapath_MV1_int_v_7__5_,
         constructing_unit_Datapath_MV1_int_v_7__6_,
         constructing_unit_Datapath_MV1_int_v_7__7_,
         constructing_unit_Datapath_MV1_int_v_7__8_,
         constructing_unit_Datapath_MV1_int_v_7__9_,
         constructing_unit_Datapath_MV1_int_v_7__10_,
         constructing_unit_Datapath_MV1_int_v_8__0_,
         constructing_unit_Datapath_MV1_int_v_8__1_,
         constructing_unit_Datapath_MV1_int_v_8__2_,
         constructing_unit_Datapath_MV1_int_v_8__3_,
         constructing_unit_Datapath_MV1_int_v_8__4_,
         constructing_unit_Datapath_MV1_int_v_8__5_,
         constructing_unit_Datapath_MV1_int_v_8__6_,
         constructing_unit_Datapath_MV1_int_v_8__7_,
         constructing_unit_Datapath_MV1_int_v_8__8_,
         constructing_unit_Datapath_MV1_int_v_8__9_,
         constructing_unit_Datapath_MV1_int_v_8__10_,
         constructing_unit_Datapath_MV1_int_v_9__0_,
         constructing_unit_Datapath_MV1_int_v_9__1_,
         constructing_unit_Datapath_MV1_int_v_9__2_,
         constructing_unit_Datapath_MV1_int_v_9__3_,
         constructing_unit_Datapath_MV1_int_v_9__4_,
         constructing_unit_Datapath_MV1_int_v_9__5_,
         constructing_unit_Datapath_MV1_int_v_9__6_,
         constructing_unit_Datapath_MV1_int_v_9__7_,
         constructing_unit_Datapath_MV1_int_v_9__8_,
         constructing_unit_Datapath_MV1_int_v_9__9_,
         constructing_unit_Datapath_MV1_int_v_9__10_,
         constructing_unit_Datapath_MV1_int_v_10__0_,
         constructing_unit_Datapath_MV1_int_v_10__1_,
         constructing_unit_Datapath_MV1_int_v_10__2_,
         constructing_unit_Datapath_MV1_int_v_10__3_,
         constructing_unit_Datapath_MV1_int_v_10__4_,
         constructing_unit_Datapath_MV1_int_v_10__5_,
         constructing_unit_Datapath_MV1_int_v_10__6_,
         constructing_unit_Datapath_MV1_int_v_10__7_,
         constructing_unit_Datapath_MV1_int_v_10__8_,
         constructing_unit_Datapath_MV1_int_v_10__9_,
         constructing_unit_Datapath_MV1_int_v_10__10_,
         constructing_unit_Datapath_MV1_int_v_11__0_,
         constructing_unit_Datapath_MV1_int_v_11__1_,
         constructing_unit_Datapath_MV1_int_v_11__2_,
         constructing_unit_Datapath_MV1_int_v_11__3_,
         constructing_unit_Datapath_MV1_int_v_11__4_,
         constructing_unit_Datapath_MV1_int_v_11__5_,
         constructing_unit_Datapath_MV1_int_v_11__6_,
         constructing_unit_Datapath_MV1_int_v_11__7_,
         constructing_unit_Datapath_MV1_int_v_11__8_,
         constructing_unit_Datapath_MV1_int_v_11__9_,
         constructing_unit_Datapath_MV1_int_v_11__10_,
         constructing_unit_Datapath_MV1_int_v_12__0_,
         constructing_unit_Datapath_MV1_int_v_12__1_,
         constructing_unit_Datapath_MV1_int_v_12__2_,
         constructing_unit_Datapath_MV1_int_v_12__3_,
         constructing_unit_Datapath_MV1_int_v_12__4_,
         constructing_unit_Datapath_MV1_int_v_12__5_,
         constructing_unit_Datapath_MV1_int_v_12__6_,
         constructing_unit_Datapath_MV1_int_v_12__7_,
         constructing_unit_Datapath_MV1_int_v_12__8_,
         constructing_unit_Datapath_MV1_int_v_12__9_,
         constructing_unit_Datapath_MV1_int_v_12__10_,
         constructing_unit_Datapath_MV1_int_v_13__0_,
         constructing_unit_Datapath_MV1_int_v_13__1_,
         constructing_unit_Datapath_MV1_int_v_13__2_,
         constructing_unit_Datapath_MV1_int_v_13__3_,
         constructing_unit_Datapath_MV1_int_v_13__4_,
         constructing_unit_Datapath_MV1_int_v_13__5_,
         constructing_unit_Datapath_MV1_int_v_13__6_,
         constructing_unit_Datapath_MV1_int_v_13__7_,
         constructing_unit_Datapath_MV1_int_v_13__8_,
         constructing_unit_Datapath_MV1_int_v_13__9_,
         constructing_unit_Datapath_MV1_int_v_13__10_,
         constructing_unit_Datapath_L_sub1_sub_19_n12,
         constructing_unit_Datapath_L_sub1_sub_19_n11,
         constructing_unit_Datapath_L_sub1_sub_19_n10,
         constructing_unit_Datapath_L_sub1_sub_19_n9,
         constructing_unit_Datapath_L_sub1_sub_19_n8,
         constructing_unit_Datapath_L_sub1_sub_19_n7,
         constructing_unit_Datapath_L_sub1_sub_19_n6,
         constructing_unit_Datapath_L_sub1_sub_19_n5,
         constructing_unit_Datapath_L_sub1_sub_19_n4,
         constructing_unit_Datapath_L_sub1_sub_19_n3,
         constructing_unit_Datapath_L_sub1_sub_19_n2,
         constructing_unit_Datapath_L_sub1_sub_19_n1,
         constructing_unit_Datapath_mv1v_mv0v_REG_0_n1,
         constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1,
         constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1,
         constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1,
         constructing_unit_Datapath_h_sample_n1,
         constructing_unit_Datapath_w_sample_n1,
         constructing_unit_Datapath_hOw_n4, constructing_unit_Datapath_hOw_n3,
         constructing_unit_Datapath_hOw_n2, constructing_unit_Datapath_hOw_n1,
         constructing_unit_Datapath_hOw_n12,
         constructing_unit_Datapath_hOw_n11,
         constructing_unit_Datapath_hOw_n10, constructing_unit_Datapath_hOw_n9,
         constructing_unit_Datapath_hOw_RSH_SH_en,
         constructing_unit_Datapath_hOw_cmd_0_,
         constructing_unit_Datapath_hOw_cmd_1_,
         constructing_unit_Datapath_hOw_FF_X_1_n1,
         constructing_unit_Datapath_hOw_FF_X_2_n1,
         constructing_unit_Datapath_hOw_FF_X_3_n1,
         constructing_unit_Datapath_hOw_cmd_RSH_n3,
         constructing_unit_Datapath_hOw_cmd_RSH_n2,
         constructing_unit_Datapath_hOw_cmd_RSH_n1,
         constructing_unit_Datapath_hOw_cmd_RSH_n8,
         constructing_unit_Datapath_hOw_cmd_RSH_n7,
         constructing_unit_Datapath_hOw_cmd_RSH_n6,
         constructing_unit_Datapath_hOw_cmd_RSH_n5,
         constructing_unit_Datapath_hOw_cmd_RSH_n4,
         constructing_unit_Datapath_hOw_RSH_n13,
         constructing_unit_Datapath_hOw_RSH_n12,
         constructing_unit_Datapath_hOw_RSH_n11,
         constructing_unit_Datapath_hOw_RSH_n10,
         constructing_unit_Datapath_hOw_RSH_n9,
         constructing_unit_Datapath_hOw_RSH_n3,
         constructing_unit_Datapath_hOw_RSH_n2,
         constructing_unit_Datapath_hOw_RSH_n1,
         constructing_unit_Datapath_L_LR_SH2_n16,
         constructing_unit_Datapath_L_LR_SH2_n15,
         constructing_unit_Datapath_L_LR_SH2_n30,
         constructing_unit_Datapath_L_LR_SH2_n29,
         constructing_unit_Datapath_L_LR_SH2_n28,
         constructing_unit_Datapath_L_LR_SH2_n27,
         constructing_unit_Datapath_L_LR_SH2_n26,
         constructing_unit_Datapath_L_LR_SH2_n25,
         constructing_unit_Datapath_L_LR_SH2_n24,
         constructing_unit_Datapath_L_LR_SH2_n23,
         constructing_unit_Datapath_L_LR_SH2_n22,
         constructing_unit_Datapath_L_LR_SH2_n21,
         constructing_unit_Datapath_L_LR_SH2_n20,
         constructing_unit_Datapath_L_LR_SH2_n19,
         constructing_unit_Datapath_L_LR_SH2_n18,
         constructing_unit_Datapath_L_LR_SH2_n17,
         constructing_unit_Datapath_L_LR_SH2_SH_en2,
         constructing_unit_Datapath_L_LR_SH2_SH_en,
         constructing_unit_Datapath_L_LR_SH2_shift_amt_int_0_,
         constructing_unit_Datapath_L_LR_SH2_shift_amt_int_1_,
         constructing_unit_Datapath_L_LR_SH2_shift_dir_int_1_,
         constructing_unit_Datapath_L_LR_SH2_shift_dir_int_2_,
         constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_,
         constructing_unit_Datapath_L_LR_SH2_FF_X_1_n1,
         constructing_unit_Datapath_L_LR_SH2_FF_X_2_n1,
         constructing_unit_Datapath_L_LR_SH2_FF_X_3_n1,
         constructing_unit_Datapath_L_LR_SH2_shift_amt_sample_n1,
         constructing_unit_Datapath_L_LR_SH2_SH_en2_sampling_n1,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n16,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n15,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n14,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n13,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n12,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n11,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n10,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n9,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n8,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n7,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n6,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n5,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n4,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n2,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n1,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n40,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n39,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n38,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n37,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n36,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n35,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n34,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n33,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n32,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n31,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n30,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n29,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n28,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n27,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n26,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n25,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n24,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n23,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n22,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n21,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n20,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n19,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n18,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n17,
         constructing_unit_Datapath_L_LR_SH2_RSH_first_n3,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n65,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n64,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n63,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n62,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n61,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n60,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n59,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n58,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n57,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n56,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n55,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n54,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n53,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n52,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n51,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n50,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n49,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n48,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n47,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n46,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n45,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n44,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n43,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n42,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n41,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n16,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n15,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n14,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n13,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n12,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n11,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n10,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n9,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n8,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n7,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n6,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n5,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n4,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n2,
         constructing_unit_Datapath_L_LR_SH2_RSH_second_n1,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n15,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n14,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n13,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n12,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n11,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n10,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n9,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n8,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n7,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n6,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n5,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n4,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n3,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n1,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n42,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n41,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n40,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n39,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n38,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n37,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n36,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n35,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n34,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n33,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n32,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n31,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n30,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n29,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n28,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n27,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n26,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n25,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n24,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n23,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n22,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n21,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n20,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n19,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n18,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n17,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n16,
         constructing_unit_Datapath_L_LR_SH2_LSH_first_n2,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n16,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n15,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n14,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n13,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n12,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n11,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n10,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n9,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n8,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n7,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n6,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n5,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n4,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n3,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n1,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n45,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n44,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n43,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n42,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n41,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n40,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n39,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n38,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n37,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n36,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n35,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n34,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n33,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n32,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n31,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n30,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n29,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n28,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n27,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n26,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n25,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n24,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n23,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n22,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n21,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n20,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n19,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n18,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n17,
         constructing_unit_Datapath_L_LR_SH2_LSH_second_n2,
         constructing_unit_Datapath_diff_mult_v_int_samp_n1,
         constructing_unit_Datapath_MV0_int_h_ext_sample_n1,
         constructing_unit_Datapath_L_sub2_sub_19_n15,
         constructing_unit_Datapath_L_sub2_sub_19_n14,
         constructing_unit_Datapath_L_sub2_sub_19_n13,
         constructing_unit_Datapath_L_sub2_sub_19_n12,
         constructing_unit_Datapath_L_sub2_sub_19_n11,
         constructing_unit_Datapath_L_sub2_sub_19_n10,
         constructing_unit_Datapath_L_sub2_sub_19_n9,
         constructing_unit_Datapath_L_sub2_sub_19_n8,
         constructing_unit_Datapath_L_sub2_sub_19_n7,
         constructing_unit_Datapath_L_sub2_sub_19_n6,
         constructing_unit_Datapath_L_sub2_sub_19_n5,
         constructing_unit_Datapath_L_sub2_sub_19_n4,
         constructing_unit_Datapath_L_sub2_sub_19_n3,
         constructing_unit_Datapath_L_sub2_sub_19_n2,
         constructing_unit_Datapath_L_sub2_sub_19_n1,
         constructing_unit_Datapath_MV2p_int_h_sample_n1,
         constructing_unit_Datapath_MV2_int_h_ext_sample_n2,
         constructing_unit_Datapath_MV2_int_h_ext_sample_n1,
         constructing_unit_Datapath_L_subD_sub_19_n16,
         constructing_unit_Datapath_L_subD_sub_19_n15,
         constructing_unit_Datapath_L_subD_sub_19_n14,
         constructing_unit_Datapath_L_subD_sub_19_n13,
         constructing_unit_Datapath_L_subD_sub_19_n12,
         constructing_unit_Datapath_L_subD_sub_19_n11,
         constructing_unit_Datapath_L_subD_sub_19_n10,
         constructing_unit_Datapath_L_subD_sub_19_n9,
         constructing_unit_Datapath_L_subD_sub_19_n8,
         constructing_unit_Datapath_L_subD_sub_19_n7,
         constructing_unit_Datapath_L_subD_sub_19_n6,
         constructing_unit_Datapath_L_subD_sub_19_n5,
         constructing_unit_Datapath_L_subD_sub_19_n4,
         constructing_unit_Datapath_L_subD_sub_19_n3,
         constructing_unit_Datapath_L_subD_sub_19_n2,
         constructing_unit_Datapath_L_subD_sub_19_n1,
         constructing_unit_Datapath_L_subD_sub_19_DIFF_15_,
         constructing_unit_Datapath_D_h_sample_n2,
         constructing_unit_Datapath_D_h_sample_n1,
         constructing_unit_Datapath_L_squarer_product_29_,
         constructing_unit_Datapath_L_squarer_mult_13_n848,
         constructing_unit_Datapath_L_squarer_mult_13_n847,
         constructing_unit_Datapath_L_squarer_mult_13_n846,
         constructing_unit_Datapath_L_squarer_mult_13_n845,
         constructing_unit_Datapath_L_squarer_mult_13_n844,
         constructing_unit_Datapath_L_squarer_mult_13_n843,
         constructing_unit_Datapath_L_squarer_mult_13_n842,
         constructing_unit_Datapath_L_squarer_mult_13_n841,
         constructing_unit_Datapath_L_squarer_mult_13_n840,
         constructing_unit_Datapath_L_squarer_mult_13_n839,
         constructing_unit_Datapath_L_squarer_mult_13_n838,
         constructing_unit_Datapath_L_squarer_mult_13_n837,
         constructing_unit_Datapath_L_squarer_mult_13_n836,
         constructing_unit_Datapath_L_squarer_mult_13_n835,
         constructing_unit_Datapath_L_squarer_mult_13_n834,
         constructing_unit_Datapath_L_squarer_mult_13_n833,
         constructing_unit_Datapath_L_squarer_mult_13_n832,
         constructing_unit_Datapath_L_squarer_mult_13_n831,
         constructing_unit_Datapath_L_squarer_mult_13_n830,
         constructing_unit_Datapath_L_squarer_mult_13_n829,
         constructing_unit_Datapath_L_squarer_mult_13_n828,
         constructing_unit_Datapath_L_squarer_mult_13_n827,
         constructing_unit_Datapath_L_squarer_mult_13_n826,
         constructing_unit_Datapath_L_squarer_mult_13_n825,
         constructing_unit_Datapath_L_squarer_mult_13_n824,
         constructing_unit_Datapath_L_squarer_mult_13_n823,
         constructing_unit_Datapath_L_squarer_mult_13_n822,
         constructing_unit_Datapath_L_squarer_mult_13_n821,
         constructing_unit_Datapath_L_squarer_mult_13_n820,
         constructing_unit_Datapath_L_squarer_mult_13_n819,
         constructing_unit_Datapath_L_squarer_mult_13_n818,
         constructing_unit_Datapath_L_squarer_mult_13_n817,
         constructing_unit_Datapath_L_squarer_mult_13_n816,
         constructing_unit_Datapath_L_squarer_mult_13_n815,
         constructing_unit_Datapath_L_squarer_mult_13_n814,
         constructing_unit_Datapath_L_squarer_mult_13_n813,
         constructing_unit_Datapath_L_squarer_mult_13_n812,
         constructing_unit_Datapath_L_squarer_mult_13_n811,
         constructing_unit_Datapath_L_squarer_mult_13_n810,
         constructing_unit_Datapath_L_squarer_mult_13_n809,
         constructing_unit_Datapath_L_squarer_mult_13_n808,
         constructing_unit_Datapath_L_squarer_mult_13_n807,
         constructing_unit_Datapath_L_squarer_mult_13_n806,
         constructing_unit_Datapath_L_squarer_mult_13_n805,
         constructing_unit_Datapath_L_squarer_mult_13_n804,
         constructing_unit_Datapath_L_squarer_mult_13_n803,
         constructing_unit_Datapath_L_squarer_mult_13_n802,
         constructing_unit_Datapath_L_squarer_mult_13_n801,
         constructing_unit_Datapath_L_squarer_mult_13_n800,
         constructing_unit_Datapath_L_squarer_mult_13_n799,
         constructing_unit_Datapath_L_squarer_mult_13_n798,
         constructing_unit_Datapath_L_squarer_mult_13_n797,
         constructing_unit_Datapath_L_squarer_mult_13_n796,
         constructing_unit_Datapath_L_squarer_mult_13_n795,
         constructing_unit_Datapath_L_squarer_mult_13_n794,
         constructing_unit_Datapath_L_squarer_mult_13_n793,
         constructing_unit_Datapath_L_squarer_mult_13_n792,
         constructing_unit_Datapath_L_squarer_mult_13_n791,
         constructing_unit_Datapath_L_squarer_mult_13_n790,
         constructing_unit_Datapath_L_squarer_mult_13_n789,
         constructing_unit_Datapath_L_squarer_mult_13_n788,
         constructing_unit_Datapath_L_squarer_mult_13_n787,
         constructing_unit_Datapath_L_squarer_mult_13_n786,
         constructing_unit_Datapath_L_squarer_mult_13_n785,
         constructing_unit_Datapath_L_squarer_mult_13_n784,
         constructing_unit_Datapath_L_squarer_mult_13_n783,
         constructing_unit_Datapath_L_squarer_mult_13_n782,
         constructing_unit_Datapath_L_squarer_mult_13_n781,
         constructing_unit_Datapath_L_squarer_mult_13_n780,
         constructing_unit_Datapath_L_squarer_mult_13_n779,
         constructing_unit_Datapath_L_squarer_mult_13_n778,
         constructing_unit_Datapath_L_squarer_mult_13_n777,
         constructing_unit_Datapath_L_squarer_mult_13_n776,
         constructing_unit_Datapath_L_squarer_mult_13_n775,
         constructing_unit_Datapath_L_squarer_mult_13_n774,
         constructing_unit_Datapath_L_squarer_mult_13_n773,
         constructing_unit_Datapath_L_squarer_mult_13_n772,
         constructing_unit_Datapath_L_squarer_mult_13_n771,
         constructing_unit_Datapath_L_squarer_mult_13_n770,
         constructing_unit_Datapath_L_squarer_mult_13_n769,
         constructing_unit_Datapath_L_squarer_mult_13_n768,
         constructing_unit_Datapath_L_squarer_mult_13_n767,
         constructing_unit_Datapath_L_squarer_mult_13_n766,
         constructing_unit_Datapath_L_squarer_mult_13_n765,
         constructing_unit_Datapath_L_squarer_mult_13_n764,
         constructing_unit_Datapath_L_squarer_mult_13_n763,
         constructing_unit_Datapath_L_squarer_mult_13_n762,
         constructing_unit_Datapath_L_squarer_mult_13_n761,
         constructing_unit_Datapath_L_squarer_mult_13_n760,
         constructing_unit_Datapath_L_squarer_mult_13_n759,
         constructing_unit_Datapath_L_squarer_mult_13_n758,
         constructing_unit_Datapath_L_squarer_mult_13_n757,
         constructing_unit_Datapath_L_squarer_mult_13_n756,
         constructing_unit_Datapath_L_squarer_mult_13_n755,
         constructing_unit_Datapath_L_squarer_mult_13_n754,
         constructing_unit_Datapath_L_squarer_mult_13_n753,
         constructing_unit_Datapath_L_squarer_mult_13_n752,
         constructing_unit_Datapath_L_squarer_mult_13_n751,
         constructing_unit_Datapath_L_squarer_mult_13_n750,
         constructing_unit_Datapath_L_squarer_mult_13_n749,
         constructing_unit_Datapath_L_squarer_mult_13_n748,
         constructing_unit_Datapath_L_squarer_mult_13_n747,
         constructing_unit_Datapath_L_squarer_mult_13_n746,
         constructing_unit_Datapath_L_squarer_mult_13_n745,
         constructing_unit_Datapath_L_squarer_mult_13_n744,
         constructing_unit_Datapath_L_squarer_mult_13_n743,
         constructing_unit_Datapath_L_squarer_mult_13_n742,
         constructing_unit_Datapath_L_squarer_mult_13_n741,
         constructing_unit_Datapath_L_squarer_mult_13_n740,
         constructing_unit_Datapath_L_squarer_mult_13_n739,
         constructing_unit_Datapath_L_squarer_mult_13_n738,
         constructing_unit_Datapath_L_squarer_mult_13_n737,
         constructing_unit_Datapath_L_squarer_mult_13_n736,
         constructing_unit_Datapath_L_squarer_mult_13_n735,
         constructing_unit_Datapath_L_squarer_mult_13_n734,
         constructing_unit_Datapath_L_squarer_mult_13_n733,
         constructing_unit_Datapath_L_squarer_mult_13_n732,
         constructing_unit_Datapath_L_squarer_mult_13_n731,
         constructing_unit_Datapath_L_squarer_mult_13_n730,
         constructing_unit_Datapath_L_squarer_mult_13_n729,
         constructing_unit_Datapath_L_squarer_mult_13_n728,
         constructing_unit_Datapath_L_squarer_mult_13_n727,
         constructing_unit_Datapath_L_squarer_mult_13_n726,
         constructing_unit_Datapath_L_squarer_mult_13_n725,
         constructing_unit_Datapath_L_squarer_mult_13_n724,
         constructing_unit_Datapath_L_squarer_mult_13_n723,
         constructing_unit_Datapath_L_squarer_mult_13_n722,
         constructing_unit_Datapath_L_squarer_mult_13_n721,
         constructing_unit_Datapath_L_squarer_mult_13_n720,
         constructing_unit_Datapath_L_squarer_mult_13_n719,
         constructing_unit_Datapath_L_squarer_mult_13_n718,
         constructing_unit_Datapath_L_squarer_mult_13_n717,
         constructing_unit_Datapath_L_squarer_mult_13_n716,
         constructing_unit_Datapath_L_squarer_mult_13_n715,
         constructing_unit_Datapath_L_squarer_mult_13_n714,
         constructing_unit_Datapath_L_squarer_mult_13_n713,
         constructing_unit_Datapath_L_squarer_mult_13_n712,
         constructing_unit_Datapath_L_squarer_mult_13_n711,
         constructing_unit_Datapath_L_squarer_mult_13_n710,
         constructing_unit_Datapath_L_squarer_mult_13_n709,
         constructing_unit_Datapath_L_squarer_mult_13_n708,
         constructing_unit_Datapath_L_squarer_mult_13_n707,
         constructing_unit_Datapath_L_squarer_mult_13_n706,
         constructing_unit_Datapath_L_squarer_mult_13_n705,
         constructing_unit_Datapath_L_squarer_mult_13_n704,
         constructing_unit_Datapath_L_squarer_mult_13_n703,
         constructing_unit_Datapath_L_squarer_mult_13_n702,
         constructing_unit_Datapath_L_squarer_mult_13_n701,
         constructing_unit_Datapath_L_squarer_mult_13_n700,
         constructing_unit_Datapath_L_squarer_mult_13_n699,
         constructing_unit_Datapath_L_squarer_mult_13_n698,
         constructing_unit_Datapath_L_squarer_mult_13_n697,
         constructing_unit_Datapath_L_squarer_mult_13_n696,
         constructing_unit_Datapath_L_squarer_mult_13_n695,
         constructing_unit_Datapath_L_squarer_mult_13_n694,
         constructing_unit_Datapath_L_squarer_mult_13_n693,
         constructing_unit_Datapath_L_squarer_mult_13_n692,
         constructing_unit_Datapath_L_squarer_mult_13_n691,
         constructing_unit_Datapath_L_squarer_mult_13_n690,
         constructing_unit_Datapath_L_squarer_mult_13_n689,
         constructing_unit_Datapath_L_squarer_mult_13_n688,
         constructing_unit_Datapath_L_squarer_mult_13_n687,
         constructing_unit_Datapath_L_squarer_mult_13_n686,
         constructing_unit_Datapath_L_squarer_mult_13_n685,
         constructing_unit_Datapath_L_squarer_mult_13_n684,
         constructing_unit_Datapath_L_squarer_mult_13_n683,
         constructing_unit_Datapath_L_squarer_mult_13_n682,
         constructing_unit_Datapath_L_squarer_mult_13_n681,
         constructing_unit_Datapath_L_squarer_mult_13_n680,
         constructing_unit_Datapath_L_squarer_mult_13_n679,
         constructing_unit_Datapath_L_squarer_mult_13_n678,
         constructing_unit_Datapath_L_squarer_mult_13_n677,
         constructing_unit_Datapath_L_squarer_mult_13_n676,
         constructing_unit_Datapath_L_squarer_mult_13_n675,
         constructing_unit_Datapath_L_squarer_mult_13_n674,
         constructing_unit_Datapath_L_squarer_mult_13_n673,
         constructing_unit_Datapath_L_squarer_mult_13_n672,
         constructing_unit_Datapath_L_squarer_mult_13_n671,
         constructing_unit_Datapath_L_squarer_mult_13_n670,
         constructing_unit_Datapath_L_squarer_mult_13_n669,
         constructing_unit_Datapath_L_squarer_mult_13_n668,
         constructing_unit_Datapath_L_squarer_mult_13_n667,
         constructing_unit_Datapath_L_squarer_mult_13_n666,
         constructing_unit_Datapath_L_squarer_mult_13_n665,
         constructing_unit_Datapath_L_squarer_mult_13_n664,
         constructing_unit_Datapath_L_squarer_mult_13_n663,
         constructing_unit_Datapath_L_squarer_mult_13_n662,
         constructing_unit_Datapath_L_squarer_mult_13_n661,
         constructing_unit_Datapath_L_squarer_mult_13_n660,
         constructing_unit_Datapath_L_squarer_mult_13_n659,
         constructing_unit_Datapath_L_squarer_mult_13_product_28_,
         constructing_unit_Datapath_L_squarer_mult_13_product_27_,
         constructing_unit_Datapath_L_squarer_mult_13_n411,
         constructing_unit_Datapath_L_squarer_mult_13_n410,
         constructing_unit_Datapath_L_squarer_mult_13_n409,
         constructing_unit_Datapath_L_squarer_mult_13_n408,
         constructing_unit_Datapath_L_squarer_mult_13_n407,
         constructing_unit_Datapath_L_squarer_mult_13_n406,
         constructing_unit_Datapath_L_squarer_mult_13_n405,
         constructing_unit_Datapath_L_squarer_mult_13_n404,
         constructing_unit_Datapath_L_squarer_mult_13_n403,
         constructing_unit_Datapath_L_squarer_mult_13_n402,
         constructing_unit_Datapath_L_squarer_mult_13_n401,
         constructing_unit_Datapath_L_squarer_mult_13_n400,
         constructing_unit_Datapath_L_squarer_mult_13_n399,
         constructing_unit_Datapath_L_squarer_mult_13_n398,
         constructing_unit_Datapath_L_squarer_mult_13_n396,
         constructing_unit_Datapath_L_squarer_mult_13_n395,
         constructing_unit_Datapath_L_squarer_mult_13_n394,
         constructing_unit_Datapath_L_squarer_mult_13_n393,
         constructing_unit_Datapath_L_squarer_mult_13_n392,
         constructing_unit_Datapath_L_squarer_mult_13_n391,
         constructing_unit_Datapath_L_squarer_mult_13_n390,
         constructing_unit_Datapath_L_squarer_mult_13_n389,
         constructing_unit_Datapath_L_squarer_mult_13_n388,
         constructing_unit_Datapath_L_squarer_mult_13_n387,
         constructing_unit_Datapath_L_squarer_mult_13_n386,
         constructing_unit_Datapath_L_squarer_mult_13_n385,
         constructing_unit_Datapath_L_squarer_mult_13_n384,
         constructing_unit_Datapath_L_squarer_mult_13_n383,
         constructing_unit_Datapath_L_squarer_mult_13_n381,
         constructing_unit_Datapath_L_squarer_mult_13_n380,
         constructing_unit_Datapath_L_squarer_mult_13_n379,
         constructing_unit_Datapath_L_squarer_mult_13_n378,
         constructing_unit_Datapath_L_squarer_mult_13_n377,
         constructing_unit_Datapath_L_squarer_mult_13_n376,
         constructing_unit_Datapath_L_squarer_mult_13_n375,
         constructing_unit_Datapath_L_squarer_mult_13_n374,
         constructing_unit_Datapath_L_squarer_mult_13_n373,
         constructing_unit_Datapath_L_squarer_mult_13_n372,
         constructing_unit_Datapath_L_squarer_mult_13_n371,
         constructing_unit_Datapath_L_squarer_mult_13_n370,
         constructing_unit_Datapath_L_squarer_mult_13_n369,
         constructing_unit_Datapath_L_squarer_mult_13_n368,
         constructing_unit_Datapath_L_squarer_mult_13_n366,
         constructing_unit_Datapath_L_squarer_mult_13_n365,
         constructing_unit_Datapath_L_squarer_mult_13_n364,
         constructing_unit_Datapath_L_squarer_mult_13_n363,
         constructing_unit_Datapath_L_squarer_mult_13_n362,
         constructing_unit_Datapath_L_squarer_mult_13_n361,
         constructing_unit_Datapath_L_squarer_mult_13_n360,
         constructing_unit_Datapath_L_squarer_mult_13_n359,
         constructing_unit_Datapath_L_squarer_mult_13_n358,
         constructing_unit_Datapath_L_squarer_mult_13_n357,
         constructing_unit_Datapath_L_squarer_mult_13_n356,
         constructing_unit_Datapath_L_squarer_mult_13_n355,
         constructing_unit_Datapath_L_squarer_mult_13_n354,
         constructing_unit_Datapath_L_squarer_mult_13_n353,
         constructing_unit_Datapath_L_squarer_mult_13_n351,
         constructing_unit_Datapath_L_squarer_mult_13_n350,
         constructing_unit_Datapath_L_squarer_mult_13_n349,
         constructing_unit_Datapath_L_squarer_mult_13_n348,
         constructing_unit_Datapath_L_squarer_mult_13_n347,
         constructing_unit_Datapath_L_squarer_mult_13_n346,
         constructing_unit_Datapath_L_squarer_mult_13_n345,
         constructing_unit_Datapath_L_squarer_mult_13_n344,
         constructing_unit_Datapath_L_squarer_mult_13_n343,
         constructing_unit_Datapath_L_squarer_mult_13_n342,
         constructing_unit_Datapath_L_squarer_mult_13_n341,
         constructing_unit_Datapath_L_squarer_mult_13_n340,
         constructing_unit_Datapath_L_squarer_mult_13_n339,
         constructing_unit_Datapath_L_squarer_mult_13_n338,
         constructing_unit_Datapath_L_squarer_mult_13_n336,
         constructing_unit_Datapath_L_squarer_mult_13_n335,
         constructing_unit_Datapath_L_squarer_mult_13_n334,
         constructing_unit_Datapath_L_squarer_mult_13_n333,
         constructing_unit_Datapath_L_squarer_mult_13_n332,
         constructing_unit_Datapath_L_squarer_mult_13_n331,
         constructing_unit_Datapath_L_squarer_mult_13_n330,
         constructing_unit_Datapath_L_squarer_mult_13_n329,
         constructing_unit_Datapath_L_squarer_mult_13_n328,
         constructing_unit_Datapath_L_squarer_mult_13_n327,
         constructing_unit_Datapath_L_squarer_mult_13_n326,
         constructing_unit_Datapath_L_squarer_mult_13_n325,
         constructing_unit_Datapath_L_squarer_mult_13_n324,
         constructing_unit_Datapath_L_squarer_mult_13_n323,
         constructing_unit_Datapath_L_squarer_mult_13_n321,
         constructing_unit_Datapath_L_squarer_mult_13_n320,
         constructing_unit_Datapath_L_squarer_mult_13_n319,
         constructing_unit_Datapath_L_squarer_mult_13_n317,
         constructing_unit_Datapath_L_squarer_mult_13_n316,
         constructing_unit_Datapath_L_squarer_mult_13_n315,
         constructing_unit_Datapath_L_squarer_mult_13_n314,
         constructing_unit_Datapath_L_squarer_mult_13_n313,
         constructing_unit_Datapath_L_squarer_mult_13_n312,
         constructing_unit_Datapath_L_squarer_mult_13_n311,
         constructing_unit_Datapath_L_squarer_mult_13_n310,
         constructing_unit_Datapath_L_squarer_mult_13_n309,
         constructing_unit_Datapath_L_squarer_mult_13_n308,
         constructing_unit_Datapath_L_squarer_mult_13_n306,
         constructing_unit_Datapath_L_squarer_mult_13_n304,
         constructing_unit_Datapath_L_squarer_mult_13_n303,
         constructing_unit_Datapath_L_squarer_mult_13_n302,
         constructing_unit_Datapath_L_squarer_mult_13_n301,
         constructing_unit_Datapath_L_squarer_mult_13_n300,
         constructing_unit_Datapath_L_squarer_mult_13_n299,
         constructing_unit_Datapath_L_squarer_mult_13_n298,
         constructing_unit_Datapath_L_squarer_mult_13_n297,
         constructing_unit_Datapath_L_squarer_mult_13_n296,
         constructing_unit_Datapath_L_squarer_mult_13_n295,
         constructing_unit_Datapath_L_squarer_mult_13_n294,
         constructing_unit_Datapath_L_squarer_mult_13_n293,
         constructing_unit_Datapath_L_squarer_mult_13_n291,
         constructing_unit_Datapath_L_squarer_mult_13_n290,
         constructing_unit_Datapath_L_squarer_mult_13_n289,
         constructing_unit_Datapath_L_squarer_mult_13_n288,
         constructing_unit_Datapath_L_squarer_mult_13_n287,
         constructing_unit_Datapath_L_squarer_mult_13_n286,
         constructing_unit_Datapath_L_squarer_mult_13_n285,
         constructing_unit_Datapath_L_squarer_mult_13_n284,
         constructing_unit_Datapath_L_squarer_mult_13_n259,
         constructing_unit_Datapath_L_squarer_mult_13_n258,
         constructing_unit_Datapath_L_squarer_mult_13_n257,
         constructing_unit_Datapath_L_squarer_mult_13_n256,
         constructing_unit_Datapath_L_squarer_mult_13_n255,
         constructing_unit_Datapath_L_squarer_mult_13_n254,
         constructing_unit_Datapath_L_squarer_mult_13_n253,
         constructing_unit_Datapath_L_squarer_mult_13_n252,
         constructing_unit_Datapath_L_squarer_mult_13_n251,
         constructing_unit_Datapath_L_squarer_mult_13_n250,
         constructing_unit_Datapath_L_squarer_mult_13_n249,
         constructing_unit_Datapath_L_squarer_mult_13_n248,
         constructing_unit_Datapath_L_squarer_mult_13_n247,
         constructing_unit_Datapath_L_squarer_mult_13_n246,
         constructing_unit_Datapath_L_squarer_mult_13_n245,
         constructing_unit_Datapath_L_squarer_mult_13_n244,
         constructing_unit_Datapath_L_squarer_mult_13_n243,
         constructing_unit_Datapath_L_squarer_mult_13_n242,
         constructing_unit_Datapath_L_squarer_mult_13_n241,
         constructing_unit_Datapath_L_squarer_mult_13_n240,
         constructing_unit_Datapath_L_squarer_mult_13_n239,
         constructing_unit_Datapath_L_squarer_mult_13_n238,
         constructing_unit_Datapath_L_squarer_mult_13_n237,
         constructing_unit_Datapath_L_squarer_mult_13_n236,
         constructing_unit_Datapath_L_squarer_mult_13_n235,
         constructing_unit_Datapath_L_squarer_mult_13_n234,
         constructing_unit_Datapath_L_squarer_mult_13_n233,
         constructing_unit_Datapath_L_squarer_mult_13_n232,
         constructing_unit_Datapath_L_squarer_mult_13_n231,
         constructing_unit_Datapath_L_squarer_mult_13_n230,
         constructing_unit_Datapath_L_squarer_mult_13_n229,
         constructing_unit_Datapath_L_squarer_mult_13_n228,
         constructing_unit_Datapath_L_squarer_mult_13_n227,
         constructing_unit_Datapath_L_squarer_mult_13_n226,
         constructing_unit_Datapath_L_squarer_mult_13_n225,
         constructing_unit_Datapath_L_squarer_mult_13_n224,
         constructing_unit_Datapath_L_squarer_mult_13_n223,
         constructing_unit_Datapath_L_squarer_mult_13_n222,
         constructing_unit_Datapath_L_squarer_mult_13_n221,
         constructing_unit_Datapath_L_squarer_mult_13_n220,
         constructing_unit_Datapath_L_squarer_mult_13_n219,
         constructing_unit_Datapath_L_squarer_mult_13_n218,
         constructing_unit_Datapath_L_squarer_mult_13_n217,
         constructing_unit_Datapath_L_squarer_mult_13_n216,
         constructing_unit_Datapath_L_squarer_mult_13_n215,
         constructing_unit_Datapath_L_squarer_mult_13_n214,
         constructing_unit_Datapath_L_squarer_mult_13_n213,
         constructing_unit_Datapath_L_squarer_mult_13_n212,
         constructing_unit_Datapath_L_squarer_mult_13_n211,
         constructing_unit_Datapath_L_squarer_mult_13_n210,
         constructing_unit_Datapath_L_squarer_mult_13_n209,
         constructing_unit_Datapath_L_squarer_mult_13_n208,
         constructing_unit_Datapath_L_squarer_mult_13_n207,
         constructing_unit_Datapath_L_squarer_mult_13_n206,
         constructing_unit_Datapath_L_squarer_mult_13_n205,
         constructing_unit_Datapath_L_squarer_mult_13_n204,
         constructing_unit_Datapath_L_squarer_mult_13_n203,
         constructing_unit_Datapath_L_squarer_mult_13_n202,
         constructing_unit_Datapath_L_squarer_mult_13_n201,
         constructing_unit_Datapath_L_squarer_mult_13_n200,
         constructing_unit_Datapath_L_squarer_mult_13_n199,
         constructing_unit_Datapath_L_squarer_mult_13_n198,
         constructing_unit_Datapath_L_squarer_mult_13_n197,
         constructing_unit_Datapath_L_squarer_mult_13_n196,
         constructing_unit_Datapath_L_squarer_mult_13_n195,
         constructing_unit_Datapath_L_squarer_mult_13_n194,
         constructing_unit_Datapath_L_squarer_mult_13_n193,
         constructing_unit_Datapath_L_squarer_mult_13_n192,
         constructing_unit_Datapath_L_squarer_mult_13_n191,
         constructing_unit_Datapath_L_squarer_mult_13_n190,
         constructing_unit_Datapath_L_squarer_mult_13_n189,
         constructing_unit_Datapath_L_squarer_mult_13_n188,
         constructing_unit_Datapath_L_squarer_mult_13_n187,
         constructing_unit_Datapath_L_squarer_mult_13_n186,
         constructing_unit_Datapath_L_squarer_mult_13_n185,
         constructing_unit_Datapath_L_squarer_mult_13_n184,
         constructing_unit_Datapath_L_squarer_mult_13_n183,
         constructing_unit_Datapath_L_squarer_mult_13_n182,
         constructing_unit_Datapath_L_squarer_mult_13_n181,
         constructing_unit_Datapath_L_squarer_mult_13_n180,
         constructing_unit_Datapath_L_squarer_mult_13_n179,
         constructing_unit_Datapath_L_squarer_mult_13_n178,
         constructing_unit_Datapath_L_squarer_mult_13_n177,
         constructing_unit_Datapath_L_squarer_mult_13_n176,
         constructing_unit_Datapath_L_squarer_mult_13_n175,
         constructing_unit_Datapath_L_squarer_mult_13_n174,
         constructing_unit_Datapath_L_squarer_mult_13_n173,
         constructing_unit_Datapath_L_squarer_mult_13_n172,
         constructing_unit_Datapath_L_squarer_mult_13_n171,
         constructing_unit_Datapath_L_squarer_mult_13_n170,
         constructing_unit_Datapath_L_squarer_mult_13_n169,
         constructing_unit_Datapath_L_squarer_mult_13_n168,
         constructing_unit_Datapath_L_squarer_mult_13_n167,
         constructing_unit_Datapath_L_squarer_mult_13_n166,
         constructing_unit_Datapath_L_squarer_mult_13_n165,
         constructing_unit_Datapath_L_squarer_mult_13_n164,
         constructing_unit_Datapath_L_squarer_mult_13_n163,
         constructing_unit_Datapath_L_squarer_mult_13_n162,
         constructing_unit_Datapath_L_squarer_mult_13_n160,
         constructing_unit_Datapath_L_squarer_mult_13_n159,
         constructing_unit_Datapath_L_squarer_mult_13_n158,
         constructing_unit_Datapath_L_squarer_mult_13_n157,
         constructing_unit_Datapath_L_squarer_mult_13_n156,
         constructing_unit_Datapath_L_squarer_mult_13_n155,
         constructing_unit_Datapath_L_squarer_mult_13_n154,
         constructing_unit_Datapath_L_squarer_mult_13_n153,
         constructing_unit_Datapath_L_squarer_mult_13_n152,
         constructing_unit_Datapath_L_squarer_mult_13_n151,
         constructing_unit_Datapath_L_squarer_mult_13_n150,
         constructing_unit_Datapath_L_squarer_mult_13_n149,
         constructing_unit_Datapath_L_squarer_mult_13_n148,
         constructing_unit_Datapath_L_squarer_mult_13_n147,
         constructing_unit_Datapath_L_squarer_mult_13_n146,
         constructing_unit_Datapath_L_squarer_mult_13_n145,
         constructing_unit_Datapath_L_squarer_mult_13_n144,
         constructing_unit_Datapath_L_squarer_mult_13_n143,
         constructing_unit_Datapath_L_squarer_mult_13_n142,
         constructing_unit_Datapath_L_squarer_mult_13_n141,
         constructing_unit_Datapath_L_squarer_mult_13_n140,
         constructing_unit_Datapath_L_squarer_mult_13_n139,
         constructing_unit_Datapath_L_squarer_mult_13_n138,
         constructing_unit_Datapath_L_squarer_mult_13_n137,
         constructing_unit_Datapath_L_squarer_mult_13_n136,
         constructing_unit_Datapath_L_squarer_mult_13_n134,
         constructing_unit_Datapath_L_squarer_mult_13_n133,
         constructing_unit_Datapath_L_squarer_mult_13_n132,
         constructing_unit_Datapath_L_squarer_mult_13_n131,
         constructing_unit_Datapath_L_squarer_mult_13_n130,
         constructing_unit_Datapath_L_squarer_mult_13_n129,
         constructing_unit_Datapath_L_squarer_mult_13_n128,
         constructing_unit_Datapath_L_squarer_mult_13_n127,
         constructing_unit_Datapath_L_squarer_mult_13_n126,
         constructing_unit_Datapath_L_squarer_mult_13_n125,
         constructing_unit_Datapath_L_squarer_mult_13_n124,
         constructing_unit_Datapath_L_squarer_mult_13_n123,
         constructing_unit_Datapath_L_squarer_mult_13_n122,
         constructing_unit_Datapath_L_squarer_mult_13_n121,
         constructing_unit_Datapath_L_squarer_mult_13_n120,
         constructing_unit_Datapath_L_squarer_mult_13_n119,
         constructing_unit_Datapath_L_squarer_mult_13_n118,
         constructing_unit_Datapath_L_squarer_mult_13_n117,
         constructing_unit_Datapath_L_squarer_mult_13_n116,
         constructing_unit_Datapath_L_squarer_mult_13_n115,
         constructing_unit_Datapath_L_squarer_mult_13_n114,
         constructing_unit_Datapath_L_squarer_mult_13_n112,
         constructing_unit_Datapath_L_squarer_mult_13_n111,
         constructing_unit_Datapath_L_squarer_mult_13_n110,
         constructing_unit_Datapath_L_squarer_mult_13_n109,
         constructing_unit_Datapath_L_squarer_mult_13_n108,
         constructing_unit_Datapath_L_squarer_mult_13_n107,
         constructing_unit_Datapath_L_squarer_mult_13_n106,
         constructing_unit_Datapath_L_squarer_mult_13_n105,
         constructing_unit_Datapath_L_squarer_mult_13_n104,
         constructing_unit_Datapath_L_squarer_mult_13_n103,
         constructing_unit_Datapath_L_squarer_mult_13_n102,
         constructing_unit_Datapath_L_squarer_mult_13_n101,
         constructing_unit_Datapath_L_squarer_mult_13_n100,
         constructing_unit_Datapath_L_squarer_mult_13_n99,
         constructing_unit_Datapath_L_squarer_mult_13_n98,
         constructing_unit_Datapath_L_squarer_mult_13_n97,
         constructing_unit_Datapath_L_squarer_mult_13_n96,
         constructing_unit_Datapath_L_squarer_mult_13_n94,
         constructing_unit_Datapath_L_squarer_mult_13_n93,
         constructing_unit_Datapath_L_squarer_mult_13_n92,
         constructing_unit_Datapath_L_squarer_mult_13_n91,
         constructing_unit_Datapath_L_squarer_mult_13_n90,
         constructing_unit_Datapath_L_squarer_mult_13_n89,
         constructing_unit_Datapath_L_squarer_mult_13_n88,
         constructing_unit_Datapath_L_squarer_mult_13_n87,
         constructing_unit_Datapath_L_squarer_mult_13_n86,
         constructing_unit_Datapath_L_squarer_mult_13_n85,
         constructing_unit_Datapath_L_squarer_mult_13_n84,
         constructing_unit_Datapath_L_squarer_mult_13_n83,
         constructing_unit_Datapath_L_squarer_mult_13_n82,
         constructing_unit_Datapath_L_squarer_mult_13_n80,
         constructing_unit_Datapath_L_squarer_mult_13_n79,
         constructing_unit_Datapath_L_squarer_mult_13_n78,
         constructing_unit_Datapath_L_squarer_mult_13_n77,
         constructing_unit_Datapath_L_squarer_mult_13_n76,
         constructing_unit_Datapath_L_squarer_mult_13_n75,
         constructing_unit_Datapath_L_squarer_mult_13_n74,
         constructing_unit_Datapath_L_squarer_mult_13_n73,
         constructing_unit_Datapath_L_squarer_mult_13_n72,
         constructing_unit_Datapath_L_squarer_mult_13_n70,
         constructing_unit_Datapath_L_squarer_mult_13_n69,
         constructing_unit_Datapath_L_squarer_mult_13_n68,
         constructing_unit_Datapath_L_squarer_mult_13_n67,
         constructing_unit_Datapath_L_squarer_mult_13_n66,
         constructing_unit_Datapath_L_squarer_mult_13_n63,
         constructing_unit_Datapath_L_squarer_mult_13_n62,
         constructing_unit_Datapath_L_squarer_mult_13_n61,
         constructing_unit_Datapath_L_squarer_mult_13_n60,
         constructing_unit_Datapath_L_squarer_mult_13_n59,
         constructing_unit_Datapath_L_squarer_mult_13_n58,
         constructing_unit_Datapath_L_squarer_mult_13_n57,
         constructing_unit_Datapath_L_squarer_mult_13_n56,
         constructing_unit_Datapath_L_squarer_mult_13_n55,
         constructing_unit_Datapath_L_squarer_mult_13_n54,
         constructing_unit_Datapath_L_squarer_mult_13_n53,
         constructing_unit_Datapath_L_squarer_mult_13_n52,
         constructing_unit_Datapath_L_squarer_mult_13_n51,
         constructing_unit_Datapath_L_squarer_mult_13_n50,
         constructing_unit_Datapath_L_squarer_mult_13_n49,
         constructing_unit_Datapath_L_squarer_mult_13_n48,
         constructing_unit_Datapath_L_squarer_mult_13_n47,
         constructing_unit_Datapath_L_squarer_mult_13_n46,
         constructing_unit_Datapath_L_squarer_mult_13_n45,
         constructing_unit_Datapath_L_squarer_mult_13_n44,
         constructing_unit_Datapath_L_squarer_mult_13_n43,
         constructing_unit_Datapath_L_squarer_mult_13_n42,
         constructing_unit_Datapath_L_squarer_mult_13_n41,
         constructing_unit_Datapath_L_squarer_mult_13_n40,
         constructing_unit_Datapath_L_squarer_mult_13_n39,
         constructing_unit_Datapath_L_squarer_mult_13_n38,
         constructing_unit_Datapath_R_sub1_sub_19_n12,
         constructing_unit_Datapath_R_sub1_sub_19_n11,
         constructing_unit_Datapath_R_sub1_sub_19_n10,
         constructing_unit_Datapath_R_sub1_sub_19_n9,
         constructing_unit_Datapath_R_sub1_sub_19_n8,
         constructing_unit_Datapath_R_sub1_sub_19_n7,
         constructing_unit_Datapath_R_sub1_sub_19_n6,
         constructing_unit_Datapath_R_sub1_sub_19_n5,
         constructing_unit_Datapath_R_sub1_sub_19_n4,
         constructing_unit_Datapath_R_sub1_sub_19_n3,
         constructing_unit_Datapath_R_sub1_sub_19_n2,
         constructing_unit_Datapath_R_sub1_sub_19_n1,
         constructing_unit_Datapath_mv1h_mv0h_REG_0_n1,
         constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1,
         constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1,
         constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1,
         constructing_unit_Datapath_R_LR_SH2_n44,
         constructing_unit_Datapath_R_LR_SH2_n43,
         constructing_unit_Datapath_R_LR_SH2_n42,
         constructing_unit_Datapath_R_LR_SH2_n41,
         constructing_unit_Datapath_R_LR_SH2_n40,
         constructing_unit_Datapath_R_LR_SH2_n39,
         constructing_unit_Datapath_R_LR_SH2_n38,
         constructing_unit_Datapath_R_LR_SH2_n37,
         constructing_unit_Datapath_R_LR_SH2_n36,
         constructing_unit_Datapath_R_LR_SH2_n35,
         constructing_unit_Datapath_R_LR_SH2_n34,
         constructing_unit_Datapath_R_LR_SH2_n33,
         constructing_unit_Datapath_R_LR_SH2_n32,
         constructing_unit_Datapath_R_LR_SH2_n31,
         constructing_unit_Datapath_R_LR_SH2_n16,
         constructing_unit_Datapath_R_LR_SH2_n15,
         constructing_unit_Datapath_R_LR_SH2_SH_en2,
         constructing_unit_Datapath_R_LR_SH2_SH_en,
         constructing_unit_Datapath_R_LR_SH2_shift_amt_int_0_,
         constructing_unit_Datapath_R_LR_SH2_shift_amt_int_1_,
         constructing_unit_Datapath_R_LR_SH2_shift_dir_int_1_,
         constructing_unit_Datapath_R_LR_SH2_shift_dir_int_2_,
         constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_,
         constructing_unit_Datapath_R_LR_SH2_FF_X_1_n1,
         constructing_unit_Datapath_R_LR_SH2_FF_X_2_n1,
         constructing_unit_Datapath_R_LR_SH2_FF_X_3_n1,
         constructing_unit_Datapath_R_LR_SH2_shift_amt_sample_n1,
         constructing_unit_Datapath_R_LR_SH2_SH_en2_sampling_n1,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n65,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n64,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n63,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n62,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n61,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n60,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n59,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n58,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n57,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n56,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n55,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n54,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n53,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n52,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n51,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n50,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n49,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n48,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n47,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n46,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n45,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n44,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n43,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n42,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n41,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n16,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n15,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n14,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n13,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n12,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n11,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n10,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n9,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n8,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n7,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n6,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n5,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n4,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n2,
         constructing_unit_Datapath_R_LR_SH2_RSH_first_n1,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n65,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n64,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n63,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n62,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n61,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n60,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n59,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n58,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n57,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n56,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n55,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n54,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n53,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n52,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n51,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n50,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n49,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n48,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n47,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n46,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n45,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n44,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n43,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n42,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n41,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n16,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n15,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n14,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n13,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n12,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n11,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n10,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n9,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n8,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n7,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n6,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n5,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n4,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n2,
         constructing_unit_Datapath_R_LR_SH2_RSH_second_n1,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n70,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n69,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n68,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n67,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n66,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n65,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n64,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n63,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n62,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n61,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n60,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n59,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n58,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n57,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n56,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n55,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n54,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n53,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n52,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n51,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n50,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n49,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n48,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n47,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n46,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n45,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n44,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n43,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n15,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n14,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n13,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n12,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n11,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n10,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n9,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n8,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n7,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n6,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n5,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n4,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n3,
         constructing_unit_Datapath_R_LR_SH2_LSH_first_n1,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n75,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n74,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n73,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n72,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n71,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n70,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n69,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n68,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n67,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n66,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n65,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n64,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n63,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n62,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n61,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n60,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n59,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n58,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n57,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n56,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n55,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n54,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n53,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n52,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n51,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n50,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n49,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n48,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n47,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n46,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n16,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n15,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n14,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n13,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n12,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n11,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n10,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n9,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n8,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n7,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n6,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n5,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n4,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n3,
         constructing_unit_Datapath_R_LR_SH2_LSH_second_n1,
         constructing_unit_Datapath_diff_mult_h_int_samp_n1,
         constructing_unit_Datapath_MV0_int_v_ext_sample_n1,
         constructing_unit_Datapath_R_sum_add_19_n1,
         constructing_unit_Datapath_MV2p_int_v_sample_n2,
         constructing_unit_Datapath_MV2p_int_v_sample_n1,
         constructing_unit_Datapath_MV2_int_v_ext_sample_n2,
         constructing_unit_Datapath_MV2_int_v_ext_sample_n1,
         constructing_unit_Datapath_R_subD_sub_19_n16,
         constructing_unit_Datapath_R_subD_sub_19_n15,
         constructing_unit_Datapath_R_subD_sub_19_n14,
         constructing_unit_Datapath_R_subD_sub_19_n13,
         constructing_unit_Datapath_R_subD_sub_19_n12,
         constructing_unit_Datapath_R_subD_sub_19_n11,
         constructing_unit_Datapath_R_subD_sub_19_n10,
         constructing_unit_Datapath_R_subD_sub_19_n9,
         constructing_unit_Datapath_R_subD_sub_19_n8,
         constructing_unit_Datapath_R_subD_sub_19_n7,
         constructing_unit_Datapath_R_subD_sub_19_n6,
         constructing_unit_Datapath_R_subD_sub_19_n5,
         constructing_unit_Datapath_R_subD_sub_19_n4,
         constructing_unit_Datapath_R_subD_sub_19_n3,
         constructing_unit_Datapath_R_subD_sub_19_n2,
         constructing_unit_Datapath_R_subD_sub_19_n1,
         constructing_unit_Datapath_R_subD_sub_19_DIFF_15_,
         constructing_unit_Datapath_D_v_sample_n2,
         constructing_unit_Datapath_D_v_sample_n1,
         constructing_unit_Datapath_R_squarer_product_29_,
         constructing_unit_Datapath_R_squarer_mult_13_n848,
         constructing_unit_Datapath_R_squarer_mult_13_n847,
         constructing_unit_Datapath_R_squarer_mult_13_n846,
         constructing_unit_Datapath_R_squarer_mult_13_n845,
         constructing_unit_Datapath_R_squarer_mult_13_n844,
         constructing_unit_Datapath_R_squarer_mult_13_n843,
         constructing_unit_Datapath_R_squarer_mult_13_n842,
         constructing_unit_Datapath_R_squarer_mult_13_n841,
         constructing_unit_Datapath_R_squarer_mult_13_n840,
         constructing_unit_Datapath_R_squarer_mult_13_n839,
         constructing_unit_Datapath_R_squarer_mult_13_n838,
         constructing_unit_Datapath_R_squarer_mult_13_n837,
         constructing_unit_Datapath_R_squarer_mult_13_n836,
         constructing_unit_Datapath_R_squarer_mult_13_n835,
         constructing_unit_Datapath_R_squarer_mult_13_n834,
         constructing_unit_Datapath_R_squarer_mult_13_n833,
         constructing_unit_Datapath_R_squarer_mult_13_n832,
         constructing_unit_Datapath_R_squarer_mult_13_n831,
         constructing_unit_Datapath_R_squarer_mult_13_n830,
         constructing_unit_Datapath_R_squarer_mult_13_n829,
         constructing_unit_Datapath_R_squarer_mult_13_n828,
         constructing_unit_Datapath_R_squarer_mult_13_n827,
         constructing_unit_Datapath_R_squarer_mult_13_n826,
         constructing_unit_Datapath_R_squarer_mult_13_n825,
         constructing_unit_Datapath_R_squarer_mult_13_n824,
         constructing_unit_Datapath_R_squarer_mult_13_n823,
         constructing_unit_Datapath_R_squarer_mult_13_n822,
         constructing_unit_Datapath_R_squarer_mult_13_n821,
         constructing_unit_Datapath_R_squarer_mult_13_n820,
         constructing_unit_Datapath_R_squarer_mult_13_n819,
         constructing_unit_Datapath_R_squarer_mult_13_n818,
         constructing_unit_Datapath_R_squarer_mult_13_n817,
         constructing_unit_Datapath_R_squarer_mult_13_n816,
         constructing_unit_Datapath_R_squarer_mult_13_n815,
         constructing_unit_Datapath_R_squarer_mult_13_n814,
         constructing_unit_Datapath_R_squarer_mult_13_n813,
         constructing_unit_Datapath_R_squarer_mult_13_n812,
         constructing_unit_Datapath_R_squarer_mult_13_n811,
         constructing_unit_Datapath_R_squarer_mult_13_n810,
         constructing_unit_Datapath_R_squarer_mult_13_n809,
         constructing_unit_Datapath_R_squarer_mult_13_n808,
         constructing_unit_Datapath_R_squarer_mult_13_n807,
         constructing_unit_Datapath_R_squarer_mult_13_n806,
         constructing_unit_Datapath_R_squarer_mult_13_n805,
         constructing_unit_Datapath_R_squarer_mult_13_n804,
         constructing_unit_Datapath_R_squarer_mult_13_n803,
         constructing_unit_Datapath_R_squarer_mult_13_n802,
         constructing_unit_Datapath_R_squarer_mult_13_n801,
         constructing_unit_Datapath_R_squarer_mult_13_n800,
         constructing_unit_Datapath_R_squarer_mult_13_n799,
         constructing_unit_Datapath_R_squarer_mult_13_n798,
         constructing_unit_Datapath_R_squarer_mult_13_n797,
         constructing_unit_Datapath_R_squarer_mult_13_n796,
         constructing_unit_Datapath_R_squarer_mult_13_n795,
         constructing_unit_Datapath_R_squarer_mult_13_n794,
         constructing_unit_Datapath_R_squarer_mult_13_n793,
         constructing_unit_Datapath_R_squarer_mult_13_n792,
         constructing_unit_Datapath_R_squarer_mult_13_n791,
         constructing_unit_Datapath_R_squarer_mult_13_n790,
         constructing_unit_Datapath_R_squarer_mult_13_n789,
         constructing_unit_Datapath_R_squarer_mult_13_n788,
         constructing_unit_Datapath_R_squarer_mult_13_n787,
         constructing_unit_Datapath_R_squarer_mult_13_n786,
         constructing_unit_Datapath_R_squarer_mult_13_n785,
         constructing_unit_Datapath_R_squarer_mult_13_n784,
         constructing_unit_Datapath_R_squarer_mult_13_n783,
         constructing_unit_Datapath_R_squarer_mult_13_n782,
         constructing_unit_Datapath_R_squarer_mult_13_n781,
         constructing_unit_Datapath_R_squarer_mult_13_n780,
         constructing_unit_Datapath_R_squarer_mult_13_n779,
         constructing_unit_Datapath_R_squarer_mult_13_n778,
         constructing_unit_Datapath_R_squarer_mult_13_n777,
         constructing_unit_Datapath_R_squarer_mult_13_n776,
         constructing_unit_Datapath_R_squarer_mult_13_n775,
         constructing_unit_Datapath_R_squarer_mult_13_n774,
         constructing_unit_Datapath_R_squarer_mult_13_n773,
         constructing_unit_Datapath_R_squarer_mult_13_n772,
         constructing_unit_Datapath_R_squarer_mult_13_n771,
         constructing_unit_Datapath_R_squarer_mult_13_n770,
         constructing_unit_Datapath_R_squarer_mult_13_n769,
         constructing_unit_Datapath_R_squarer_mult_13_n768,
         constructing_unit_Datapath_R_squarer_mult_13_n767,
         constructing_unit_Datapath_R_squarer_mult_13_n766,
         constructing_unit_Datapath_R_squarer_mult_13_n765,
         constructing_unit_Datapath_R_squarer_mult_13_n764,
         constructing_unit_Datapath_R_squarer_mult_13_n763,
         constructing_unit_Datapath_R_squarer_mult_13_n762,
         constructing_unit_Datapath_R_squarer_mult_13_n761,
         constructing_unit_Datapath_R_squarer_mult_13_n760,
         constructing_unit_Datapath_R_squarer_mult_13_n759,
         constructing_unit_Datapath_R_squarer_mult_13_n758,
         constructing_unit_Datapath_R_squarer_mult_13_n757,
         constructing_unit_Datapath_R_squarer_mult_13_n756,
         constructing_unit_Datapath_R_squarer_mult_13_n755,
         constructing_unit_Datapath_R_squarer_mult_13_n754,
         constructing_unit_Datapath_R_squarer_mult_13_n753,
         constructing_unit_Datapath_R_squarer_mult_13_n752,
         constructing_unit_Datapath_R_squarer_mult_13_n751,
         constructing_unit_Datapath_R_squarer_mult_13_n750,
         constructing_unit_Datapath_R_squarer_mult_13_n749,
         constructing_unit_Datapath_R_squarer_mult_13_n748,
         constructing_unit_Datapath_R_squarer_mult_13_n747,
         constructing_unit_Datapath_R_squarer_mult_13_n746,
         constructing_unit_Datapath_R_squarer_mult_13_n745,
         constructing_unit_Datapath_R_squarer_mult_13_n744,
         constructing_unit_Datapath_R_squarer_mult_13_n743,
         constructing_unit_Datapath_R_squarer_mult_13_n742,
         constructing_unit_Datapath_R_squarer_mult_13_n741,
         constructing_unit_Datapath_R_squarer_mult_13_n740,
         constructing_unit_Datapath_R_squarer_mult_13_n739,
         constructing_unit_Datapath_R_squarer_mult_13_n738,
         constructing_unit_Datapath_R_squarer_mult_13_n737,
         constructing_unit_Datapath_R_squarer_mult_13_n736,
         constructing_unit_Datapath_R_squarer_mult_13_n735,
         constructing_unit_Datapath_R_squarer_mult_13_n734,
         constructing_unit_Datapath_R_squarer_mult_13_n733,
         constructing_unit_Datapath_R_squarer_mult_13_n732,
         constructing_unit_Datapath_R_squarer_mult_13_n731,
         constructing_unit_Datapath_R_squarer_mult_13_n730,
         constructing_unit_Datapath_R_squarer_mult_13_n729,
         constructing_unit_Datapath_R_squarer_mult_13_n728,
         constructing_unit_Datapath_R_squarer_mult_13_n727,
         constructing_unit_Datapath_R_squarer_mult_13_n726,
         constructing_unit_Datapath_R_squarer_mult_13_n725,
         constructing_unit_Datapath_R_squarer_mult_13_n724,
         constructing_unit_Datapath_R_squarer_mult_13_n723,
         constructing_unit_Datapath_R_squarer_mult_13_n722,
         constructing_unit_Datapath_R_squarer_mult_13_n721,
         constructing_unit_Datapath_R_squarer_mult_13_n720,
         constructing_unit_Datapath_R_squarer_mult_13_n719,
         constructing_unit_Datapath_R_squarer_mult_13_n718,
         constructing_unit_Datapath_R_squarer_mult_13_n717,
         constructing_unit_Datapath_R_squarer_mult_13_n716,
         constructing_unit_Datapath_R_squarer_mult_13_n715,
         constructing_unit_Datapath_R_squarer_mult_13_n714,
         constructing_unit_Datapath_R_squarer_mult_13_n713,
         constructing_unit_Datapath_R_squarer_mult_13_n712,
         constructing_unit_Datapath_R_squarer_mult_13_n711,
         constructing_unit_Datapath_R_squarer_mult_13_n710,
         constructing_unit_Datapath_R_squarer_mult_13_n709,
         constructing_unit_Datapath_R_squarer_mult_13_n708,
         constructing_unit_Datapath_R_squarer_mult_13_n707,
         constructing_unit_Datapath_R_squarer_mult_13_n706,
         constructing_unit_Datapath_R_squarer_mult_13_n705,
         constructing_unit_Datapath_R_squarer_mult_13_n704,
         constructing_unit_Datapath_R_squarer_mult_13_n703,
         constructing_unit_Datapath_R_squarer_mult_13_n702,
         constructing_unit_Datapath_R_squarer_mult_13_n701,
         constructing_unit_Datapath_R_squarer_mult_13_n700,
         constructing_unit_Datapath_R_squarer_mult_13_n699,
         constructing_unit_Datapath_R_squarer_mult_13_n698,
         constructing_unit_Datapath_R_squarer_mult_13_n697,
         constructing_unit_Datapath_R_squarer_mult_13_n696,
         constructing_unit_Datapath_R_squarer_mult_13_n695,
         constructing_unit_Datapath_R_squarer_mult_13_n694,
         constructing_unit_Datapath_R_squarer_mult_13_n693,
         constructing_unit_Datapath_R_squarer_mult_13_n692,
         constructing_unit_Datapath_R_squarer_mult_13_n691,
         constructing_unit_Datapath_R_squarer_mult_13_n690,
         constructing_unit_Datapath_R_squarer_mult_13_n689,
         constructing_unit_Datapath_R_squarer_mult_13_n688,
         constructing_unit_Datapath_R_squarer_mult_13_n687,
         constructing_unit_Datapath_R_squarer_mult_13_n686,
         constructing_unit_Datapath_R_squarer_mult_13_n685,
         constructing_unit_Datapath_R_squarer_mult_13_n684,
         constructing_unit_Datapath_R_squarer_mult_13_n683,
         constructing_unit_Datapath_R_squarer_mult_13_n682,
         constructing_unit_Datapath_R_squarer_mult_13_n681,
         constructing_unit_Datapath_R_squarer_mult_13_n680,
         constructing_unit_Datapath_R_squarer_mult_13_n679,
         constructing_unit_Datapath_R_squarer_mult_13_n678,
         constructing_unit_Datapath_R_squarer_mult_13_n677,
         constructing_unit_Datapath_R_squarer_mult_13_n676,
         constructing_unit_Datapath_R_squarer_mult_13_n675,
         constructing_unit_Datapath_R_squarer_mult_13_n674,
         constructing_unit_Datapath_R_squarer_mult_13_n673,
         constructing_unit_Datapath_R_squarer_mult_13_n672,
         constructing_unit_Datapath_R_squarer_mult_13_n671,
         constructing_unit_Datapath_R_squarer_mult_13_n670,
         constructing_unit_Datapath_R_squarer_mult_13_n669,
         constructing_unit_Datapath_R_squarer_mult_13_n668,
         constructing_unit_Datapath_R_squarer_mult_13_n667,
         constructing_unit_Datapath_R_squarer_mult_13_n666,
         constructing_unit_Datapath_R_squarer_mult_13_n665,
         constructing_unit_Datapath_R_squarer_mult_13_n664,
         constructing_unit_Datapath_R_squarer_mult_13_n663,
         constructing_unit_Datapath_R_squarer_mult_13_n662,
         constructing_unit_Datapath_R_squarer_mult_13_n661,
         constructing_unit_Datapath_R_squarer_mult_13_n660,
         constructing_unit_Datapath_R_squarer_mult_13_n659,
         constructing_unit_Datapath_R_squarer_mult_13_product_28_,
         constructing_unit_Datapath_R_squarer_mult_13_product_27_,
         constructing_unit_Datapath_R_squarer_mult_13_n411,
         constructing_unit_Datapath_R_squarer_mult_13_n410,
         constructing_unit_Datapath_R_squarer_mult_13_n409,
         constructing_unit_Datapath_R_squarer_mult_13_n408,
         constructing_unit_Datapath_R_squarer_mult_13_n407,
         constructing_unit_Datapath_R_squarer_mult_13_n406,
         constructing_unit_Datapath_R_squarer_mult_13_n405,
         constructing_unit_Datapath_R_squarer_mult_13_n404,
         constructing_unit_Datapath_R_squarer_mult_13_n403,
         constructing_unit_Datapath_R_squarer_mult_13_n402,
         constructing_unit_Datapath_R_squarer_mult_13_n401,
         constructing_unit_Datapath_R_squarer_mult_13_n400,
         constructing_unit_Datapath_R_squarer_mult_13_n399,
         constructing_unit_Datapath_R_squarer_mult_13_n398,
         constructing_unit_Datapath_R_squarer_mult_13_n396,
         constructing_unit_Datapath_R_squarer_mult_13_n395,
         constructing_unit_Datapath_R_squarer_mult_13_n394,
         constructing_unit_Datapath_R_squarer_mult_13_n393,
         constructing_unit_Datapath_R_squarer_mult_13_n392,
         constructing_unit_Datapath_R_squarer_mult_13_n391,
         constructing_unit_Datapath_R_squarer_mult_13_n390,
         constructing_unit_Datapath_R_squarer_mult_13_n389,
         constructing_unit_Datapath_R_squarer_mult_13_n388,
         constructing_unit_Datapath_R_squarer_mult_13_n387,
         constructing_unit_Datapath_R_squarer_mult_13_n386,
         constructing_unit_Datapath_R_squarer_mult_13_n385,
         constructing_unit_Datapath_R_squarer_mult_13_n384,
         constructing_unit_Datapath_R_squarer_mult_13_n383,
         constructing_unit_Datapath_R_squarer_mult_13_n381,
         constructing_unit_Datapath_R_squarer_mult_13_n380,
         constructing_unit_Datapath_R_squarer_mult_13_n379,
         constructing_unit_Datapath_R_squarer_mult_13_n378,
         constructing_unit_Datapath_R_squarer_mult_13_n377,
         constructing_unit_Datapath_R_squarer_mult_13_n376,
         constructing_unit_Datapath_R_squarer_mult_13_n375,
         constructing_unit_Datapath_R_squarer_mult_13_n374,
         constructing_unit_Datapath_R_squarer_mult_13_n373,
         constructing_unit_Datapath_R_squarer_mult_13_n372,
         constructing_unit_Datapath_R_squarer_mult_13_n371,
         constructing_unit_Datapath_R_squarer_mult_13_n370,
         constructing_unit_Datapath_R_squarer_mult_13_n369,
         constructing_unit_Datapath_R_squarer_mult_13_n368,
         constructing_unit_Datapath_R_squarer_mult_13_n366,
         constructing_unit_Datapath_R_squarer_mult_13_n365,
         constructing_unit_Datapath_R_squarer_mult_13_n364,
         constructing_unit_Datapath_R_squarer_mult_13_n363,
         constructing_unit_Datapath_R_squarer_mult_13_n362,
         constructing_unit_Datapath_R_squarer_mult_13_n361,
         constructing_unit_Datapath_R_squarer_mult_13_n360,
         constructing_unit_Datapath_R_squarer_mult_13_n359,
         constructing_unit_Datapath_R_squarer_mult_13_n358,
         constructing_unit_Datapath_R_squarer_mult_13_n357,
         constructing_unit_Datapath_R_squarer_mult_13_n356,
         constructing_unit_Datapath_R_squarer_mult_13_n355,
         constructing_unit_Datapath_R_squarer_mult_13_n354,
         constructing_unit_Datapath_R_squarer_mult_13_n353,
         constructing_unit_Datapath_R_squarer_mult_13_n351,
         constructing_unit_Datapath_R_squarer_mult_13_n350,
         constructing_unit_Datapath_R_squarer_mult_13_n349,
         constructing_unit_Datapath_R_squarer_mult_13_n348,
         constructing_unit_Datapath_R_squarer_mult_13_n347,
         constructing_unit_Datapath_R_squarer_mult_13_n346,
         constructing_unit_Datapath_R_squarer_mult_13_n345,
         constructing_unit_Datapath_R_squarer_mult_13_n344,
         constructing_unit_Datapath_R_squarer_mult_13_n343,
         constructing_unit_Datapath_R_squarer_mult_13_n342,
         constructing_unit_Datapath_R_squarer_mult_13_n341,
         constructing_unit_Datapath_R_squarer_mult_13_n340,
         constructing_unit_Datapath_R_squarer_mult_13_n339,
         constructing_unit_Datapath_R_squarer_mult_13_n338,
         constructing_unit_Datapath_R_squarer_mult_13_n336,
         constructing_unit_Datapath_R_squarer_mult_13_n335,
         constructing_unit_Datapath_R_squarer_mult_13_n334,
         constructing_unit_Datapath_R_squarer_mult_13_n333,
         constructing_unit_Datapath_R_squarer_mult_13_n332,
         constructing_unit_Datapath_R_squarer_mult_13_n331,
         constructing_unit_Datapath_R_squarer_mult_13_n330,
         constructing_unit_Datapath_R_squarer_mult_13_n329,
         constructing_unit_Datapath_R_squarer_mult_13_n328,
         constructing_unit_Datapath_R_squarer_mult_13_n327,
         constructing_unit_Datapath_R_squarer_mult_13_n326,
         constructing_unit_Datapath_R_squarer_mult_13_n325,
         constructing_unit_Datapath_R_squarer_mult_13_n324,
         constructing_unit_Datapath_R_squarer_mult_13_n323,
         constructing_unit_Datapath_R_squarer_mult_13_n321,
         constructing_unit_Datapath_R_squarer_mult_13_n320,
         constructing_unit_Datapath_R_squarer_mult_13_n319,
         constructing_unit_Datapath_R_squarer_mult_13_n317,
         constructing_unit_Datapath_R_squarer_mult_13_n316,
         constructing_unit_Datapath_R_squarer_mult_13_n315,
         constructing_unit_Datapath_R_squarer_mult_13_n314,
         constructing_unit_Datapath_R_squarer_mult_13_n313,
         constructing_unit_Datapath_R_squarer_mult_13_n312,
         constructing_unit_Datapath_R_squarer_mult_13_n311,
         constructing_unit_Datapath_R_squarer_mult_13_n310,
         constructing_unit_Datapath_R_squarer_mult_13_n309,
         constructing_unit_Datapath_R_squarer_mult_13_n308,
         constructing_unit_Datapath_R_squarer_mult_13_n306,
         constructing_unit_Datapath_R_squarer_mult_13_n304,
         constructing_unit_Datapath_R_squarer_mult_13_n303,
         constructing_unit_Datapath_R_squarer_mult_13_n302,
         constructing_unit_Datapath_R_squarer_mult_13_n301,
         constructing_unit_Datapath_R_squarer_mult_13_n300,
         constructing_unit_Datapath_R_squarer_mult_13_n299,
         constructing_unit_Datapath_R_squarer_mult_13_n298,
         constructing_unit_Datapath_R_squarer_mult_13_n297,
         constructing_unit_Datapath_R_squarer_mult_13_n296,
         constructing_unit_Datapath_R_squarer_mult_13_n295,
         constructing_unit_Datapath_R_squarer_mult_13_n294,
         constructing_unit_Datapath_R_squarer_mult_13_n293,
         constructing_unit_Datapath_R_squarer_mult_13_n291,
         constructing_unit_Datapath_R_squarer_mult_13_n290,
         constructing_unit_Datapath_R_squarer_mult_13_n289,
         constructing_unit_Datapath_R_squarer_mult_13_n288,
         constructing_unit_Datapath_R_squarer_mult_13_n287,
         constructing_unit_Datapath_R_squarer_mult_13_n286,
         constructing_unit_Datapath_R_squarer_mult_13_n285,
         constructing_unit_Datapath_R_squarer_mult_13_n284,
         constructing_unit_Datapath_R_squarer_mult_13_n259,
         constructing_unit_Datapath_R_squarer_mult_13_n258,
         constructing_unit_Datapath_R_squarer_mult_13_n257,
         constructing_unit_Datapath_R_squarer_mult_13_n256,
         constructing_unit_Datapath_R_squarer_mult_13_n255,
         constructing_unit_Datapath_R_squarer_mult_13_n254,
         constructing_unit_Datapath_R_squarer_mult_13_n253,
         constructing_unit_Datapath_R_squarer_mult_13_n252,
         constructing_unit_Datapath_R_squarer_mult_13_n251,
         constructing_unit_Datapath_R_squarer_mult_13_n250,
         constructing_unit_Datapath_R_squarer_mult_13_n249,
         constructing_unit_Datapath_R_squarer_mult_13_n248,
         constructing_unit_Datapath_R_squarer_mult_13_n247,
         constructing_unit_Datapath_R_squarer_mult_13_n246,
         constructing_unit_Datapath_R_squarer_mult_13_n245,
         constructing_unit_Datapath_R_squarer_mult_13_n244,
         constructing_unit_Datapath_R_squarer_mult_13_n243,
         constructing_unit_Datapath_R_squarer_mult_13_n242,
         constructing_unit_Datapath_R_squarer_mult_13_n241,
         constructing_unit_Datapath_R_squarer_mult_13_n240,
         constructing_unit_Datapath_R_squarer_mult_13_n239,
         constructing_unit_Datapath_R_squarer_mult_13_n238,
         constructing_unit_Datapath_R_squarer_mult_13_n237,
         constructing_unit_Datapath_R_squarer_mult_13_n236,
         constructing_unit_Datapath_R_squarer_mult_13_n235,
         constructing_unit_Datapath_R_squarer_mult_13_n234,
         constructing_unit_Datapath_R_squarer_mult_13_n233,
         constructing_unit_Datapath_R_squarer_mult_13_n232,
         constructing_unit_Datapath_R_squarer_mult_13_n231,
         constructing_unit_Datapath_R_squarer_mult_13_n230,
         constructing_unit_Datapath_R_squarer_mult_13_n229,
         constructing_unit_Datapath_R_squarer_mult_13_n228,
         constructing_unit_Datapath_R_squarer_mult_13_n227,
         constructing_unit_Datapath_R_squarer_mult_13_n226,
         constructing_unit_Datapath_R_squarer_mult_13_n225,
         constructing_unit_Datapath_R_squarer_mult_13_n224,
         constructing_unit_Datapath_R_squarer_mult_13_n223,
         constructing_unit_Datapath_R_squarer_mult_13_n222,
         constructing_unit_Datapath_R_squarer_mult_13_n221,
         constructing_unit_Datapath_R_squarer_mult_13_n220,
         constructing_unit_Datapath_R_squarer_mult_13_n219,
         constructing_unit_Datapath_R_squarer_mult_13_n218,
         constructing_unit_Datapath_R_squarer_mult_13_n217,
         constructing_unit_Datapath_R_squarer_mult_13_n216,
         constructing_unit_Datapath_R_squarer_mult_13_n215,
         constructing_unit_Datapath_R_squarer_mult_13_n214,
         constructing_unit_Datapath_R_squarer_mult_13_n213,
         constructing_unit_Datapath_R_squarer_mult_13_n212,
         constructing_unit_Datapath_R_squarer_mult_13_n211,
         constructing_unit_Datapath_R_squarer_mult_13_n210,
         constructing_unit_Datapath_R_squarer_mult_13_n209,
         constructing_unit_Datapath_R_squarer_mult_13_n208,
         constructing_unit_Datapath_R_squarer_mult_13_n207,
         constructing_unit_Datapath_R_squarer_mult_13_n206,
         constructing_unit_Datapath_R_squarer_mult_13_n205,
         constructing_unit_Datapath_R_squarer_mult_13_n204,
         constructing_unit_Datapath_R_squarer_mult_13_n203,
         constructing_unit_Datapath_R_squarer_mult_13_n202,
         constructing_unit_Datapath_R_squarer_mult_13_n201,
         constructing_unit_Datapath_R_squarer_mult_13_n200,
         constructing_unit_Datapath_R_squarer_mult_13_n199,
         constructing_unit_Datapath_R_squarer_mult_13_n198,
         constructing_unit_Datapath_R_squarer_mult_13_n197,
         constructing_unit_Datapath_R_squarer_mult_13_n196,
         constructing_unit_Datapath_R_squarer_mult_13_n195,
         constructing_unit_Datapath_R_squarer_mult_13_n194,
         constructing_unit_Datapath_R_squarer_mult_13_n193,
         constructing_unit_Datapath_R_squarer_mult_13_n192,
         constructing_unit_Datapath_R_squarer_mult_13_n191,
         constructing_unit_Datapath_R_squarer_mult_13_n190,
         constructing_unit_Datapath_R_squarer_mult_13_n189,
         constructing_unit_Datapath_R_squarer_mult_13_n188,
         constructing_unit_Datapath_R_squarer_mult_13_n187,
         constructing_unit_Datapath_R_squarer_mult_13_n186,
         constructing_unit_Datapath_R_squarer_mult_13_n185,
         constructing_unit_Datapath_R_squarer_mult_13_n184,
         constructing_unit_Datapath_R_squarer_mult_13_n183,
         constructing_unit_Datapath_R_squarer_mult_13_n182,
         constructing_unit_Datapath_R_squarer_mult_13_n181,
         constructing_unit_Datapath_R_squarer_mult_13_n180,
         constructing_unit_Datapath_R_squarer_mult_13_n179,
         constructing_unit_Datapath_R_squarer_mult_13_n178,
         constructing_unit_Datapath_R_squarer_mult_13_n177,
         constructing_unit_Datapath_R_squarer_mult_13_n176,
         constructing_unit_Datapath_R_squarer_mult_13_n175,
         constructing_unit_Datapath_R_squarer_mult_13_n174,
         constructing_unit_Datapath_R_squarer_mult_13_n173,
         constructing_unit_Datapath_R_squarer_mult_13_n172,
         constructing_unit_Datapath_R_squarer_mult_13_n171,
         constructing_unit_Datapath_R_squarer_mult_13_n170,
         constructing_unit_Datapath_R_squarer_mult_13_n169,
         constructing_unit_Datapath_R_squarer_mult_13_n168,
         constructing_unit_Datapath_R_squarer_mult_13_n167,
         constructing_unit_Datapath_R_squarer_mult_13_n166,
         constructing_unit_Datapath_R_squarer_mult_13_n165,
         constructing_unit_Datapath_R_squarer_mult_13_n164,
         constructing_unit_Datapath_R_squarer_mult_13_n163,
         constructing_unit_Datapath_R_squarer_mult_13_n162,
         constructing_unit_Datapath_R_squarer_mult_13_n160,
         constructing_unit_Datapath_R_squarer_mult_13_n159,
         constructing_unit_Datapath_R_squarer_mult_13_n158,
         constructing_unit_Datapath_R_squarer_mult_13_n157,
         constructing_unit_Datapath_R_squarer_mult_13_n156,
         constructing_unit_Datapath_R_squarer_mult_13_n155,
         constructing_unit_Datapath_R_squarer_mult_13_n154,
         constructing_unit_Datapath_R_squarer_mult_13_n153,
         constructing_unit_Datapath_R_squarer_mult_13_n152,
         constructing_unit_Datapath_R_squarer_mult_13_n151,
         constructing_unit_Datapath_R_squarer_mult_13_n150,
         constructing_unit_Datapath_R_squarer_mult_13_n149,
         constructing_unit_Datapath_R_squarer_mult_13_n148,
         constructing_unit_Datapath_R_squarer_mult_13_n147,
         constructing_unit_Datapath_R_squarer_mult_13_n146,
         constructing_unit_Datapath_R_squarer_mult_13_n145,
         constructing_unit_Datapath_R_squarer_mult_13_n144,
         constructing_unit_Datapath_R_squarer_mult_13_n143,
         constructing_unit_Datapath_R_squarer_mult_13_n142,
         constructing_unit_Datapath_R_squarer_mult_13_n141,
         constructing_unit_Datapath_R_squarer_mult_13_n140,
         constructing_unit_Datapath_R_squarer_mult_13_n139,
         constructing_unit_Datapath_R_squarer_mult_13_n138,
         constructing_unit_Datapath_R_squarer_mult_13_n137,
         constructing_unit_Datapath_R_squarer_mult_13_n136,
         constructing_unit_Datapath_R_squarer_mult_13_n134,
         constructing_unit_Datapath_R_squarer_mult_13_n133,
         constructing_unit_Datapath_R_squarer_mult_13_n132,
         constructing_unit_Datapath_R_squarer_mult_13_n131,
         constructing_unit_Datapath_R_squarer_mult_13_n130,
         constructing_unit_Datapath_R_squarer_mult_13_n129,
         constructing_unit_Datapath_R_squarer_mult_13_n128,
         constructing_unit_Datapath_R_squarer_mult_13_n127,
         constructing_unit_Datapath_R_squarer_mult_13_n126,
         constructing_unit_Datapath_R_squarer_mult_13_n125,
         constructing_unit_Datapath_R_squarer_mult_13_n124,
         constructing_unit_Datapath_R_squarer_mult_13_n123,
         constructing_unit_Datapath_R_squarer_mult_13_n122,
         constructing_unit_Datapath_R_squarer_mult_13_n121,
         constructing_unit_Datapath_R_squarer_mult_13_n120,
         constructing_unit_Datapath_R_squarer_mult_13_n119,
         constructing_unit_Datapath_R_squarer_mult_13_n118,
         constructing_unit_Datapath_R_squarer_mult_13_n117,
         constructing_unit_Datapath_R_squarer_mult_13_n116,
         constructing_unit_Datapath_R_squarer_mult_13_n115,
         constructing_unit_Datapath_R_squarer_mult_13_n114,
         constructing_unit_Datapath_R_squarer_mult_13_n112,
         constructing_unit_Datapath_R_squarer_mult_13_n111,
         constructing_unit_Datapath_R_squarer_mult_13_n110,
         constructing_unit_Datapath_R_squarer_mult_13_n109,
         constructing_unit_Datapath_R_squarer_mult_13_n108,
         constructing_unit_Datapath_R_squarer_mult_13_n107,
         constructing_unit_Datapath_R_squarer_mult_13_n106,
         constructing_unit_Datapath_R_squarer_mult_13_n105,
         constructing_unit_Datapath_R_squarer_mult_13_n104,
         constructing_unit_Datapath_R_squarer_mult_13_n103,
         constructing_unit_Datapath_R_squarer_mult_13_n102,
         constructing_unit_Datapath_R_squarer_mult_13_n101,
         constructing_unit_Datapath_R_squarer_mult_13_n100,
         constructing_unit_Datapath_R_squarer_mult_13_n99,
         constructing_unit_Datapath_R_squarer_mult_13_n98,
         constructing_unit_Datapath_R_squarer_mult_13_n97,
         constructing_unit_Datapath_R_squarer_mult_13_n96,
         constructing_unit_Datapath_R_squarer_mult_13_n94,
         constructing_unit_Datapath_R_squarer_mult_13_n93,
         constructing_unit_Datapath_R_squarer_mult_13_n92,
         constructing_unit_Datapath_R_squarer_mult_13_n91,
         constructing_unit_Datapath_R_squarer_mult_13_n90,
         constructing_unit_Datapath_R_squarer_mult_13_n89,
         constructing_unit_Datapath_R_squarer_mult_13_n88,
         constructing_unit_Datapath_R_squarer_mult_13_n87,
         constructing_unit_Datapath_R_squarer_mult_13_n86,
         constructing_unit_Datapath_R_squarer_mult_13_n85,
         constructing_unit_Datapath_R_squarer_mult_13_n84,
         constructing_unit_Datapath_R_squarer_mult_13_n83,
         constructing_unit_Datapath_R_squarer_mult_13_n82,
         constructing_unit_Datapath_R_squarer_mult_13_n80,
         constructing_unit_Datapath_R_squarer_mult_13_n79,
         constructing_unit_Datapath_R_squarer_mult_13_n78,
         constructing_unit_Datapath_R_squarer_mult_13_n77,
         constructing_unit_Datapath_R_squarer_mult_13_n76,
         constructing_unit_Datapath_R_squarer_mult_13_n75,
         constructing_unit_Datapath_R_squarer_mult_13_n74,
         constructing_unit_Datapath_R_squarer_mult_13_n73,
         constructing_unit_Datapath_R_squarer_mult_13_n72,
         constructing_unit_Datapath_R_squarer_mult_13_n70,
         constructing_unit_Datapath_R_squarer_mult_13_n69,
         constructing_unit_Datapath_R_squarer_mult_13_n68,
         constructing_unit_Datapath_R_squarer_mult_13_n67,
         constructing_unit_Datapath_R_squarer_mult_13_n66,
         constructing_unit_Datapath_R_squarer_mult_13_n63,
         constructing_unit_Datapath_R_squarer_mult_13_n62,
         constructing_unit_Datapath_R_squarer_mult_13_n61,
         constructing_unit_Datapath_R_squarer_mult_13_n60,
         constructing_unit_Datapath_R_squarer_mult_13_n59,
         constructing_unit_Datapath_R_squarer_mult_13_n58,
         constructing_unit_Datapath_R_squarer_mult_13_n57,
         constructing_unit_Datapath_R_squarer_mult_13_n56,
         constructing_unit_Datapath_R_squarer_mult_13_n55,
         constructing_unit_Datapath_R_squarer_mult_13_n54,
         constructing_unit_Datapath_R_squarer_mult_13_n53,
         constructing_unit_Datapath_R_squarer_mult_13_n52,
         constructing_unit_Datapath_R_squarer_mult_13_n51,
         constructing_unit_Datapath_R_squarer_mult_13_n50,
         constructing_unit_Datapath_R_squarer_mult_13_n49,
         constructing_unit_Datapath_R_squarer_mult_13_n48,
         constructing_unit_Datapath_R_squarer_mult_13_n47,
         constructing_unit_Datapath_R_squarer_mult_13_n46,
         constructing_unit_Datapath_R_squarer_mult_13_n45,
         constructing_unit_Datapath_R_squarer_mult_13_n44,
         constructing_unit_Datapath_R_squarer_mult_13_n43,
         constructing_unit_Datapath_R_squarer_mult_13_n42,
         constructing_unit_Datapath_R_squarer_mult_13_n41,
         constructing_unit_Datapath_R_squarer_mult_13_n40,
         constructing_unit_Datapath_R_squarer_mult_13_n39,
         constructing_unit_Datapath_R_squarer_mult_13_n38,
         constructing_unit_Datapath_MV0_check_n2,
         constructing_unit_Datapath_MV0_check_n1,
         constructing_unit_Datapath_MV0_check_n10,
         constructing_unit_Datapath_MV0_check_n9,
         constructing_unit_Datapath_MV0_check_n8,
         constructing_unit_Datapath_MV0_check_n7,
         constructing_unit_Datapath_MV0_check_n6,
         constructing_unit_Datapath_MV0_check_n5,
         constructing_unit_Datapath_MV0_check_n4,
         constructing_unit_Datapath_MV0_check_n3,
         constructing_unit_Datapath_MV1_check_n18,
         constructing_unit_Datapath_MV1_check_n17,
         constructing_unit_Datapath_MV1_check_n16,
         constructing_unit_Datapath_MV1_check_n15,
         constructing_unit_Datapath_MV1_check_n14,
         constructing_unit_Datapath_MV1_check_n13,
         constructing_unit_Datapath_MV1_check_n12,
         constructing_unit_Datapath_MV1_check_n11,
         constructing_unit_Datapath_MV1_check_n2,
         constructing_unit_Datapath_MV1_check_n1,
         constructing_unit_Datapath_MV2_check_n18,
         constructing_unit_Datapath_MV2_check_n17,
         constructing_unit_Datapath_MV2_check_n16,
         constructing_unit_Datapath_MV2_check_n15,
         constructing_unit_Datapath_MV2_check_n14,
         constructing_unit_Datapath_MV2_check_n13,
         constructing_unit_Datapath_MV2_check_n12,
         constructing_unit_Datapath_MV2_check_n11,
         constructing_unit_Datapath_MV2_check_n2,
         constructing_unit_Datapath_MV2_check_n1,
         constructing_unit_Datapath_UA_flag_1st_delay_n1,
         constructing_unit_Datapath_UA_flag_delay_FFX_2_n1,
         constructing_unit_Datapath_UA_flag_delay_FFX_3_n1,
         constructing_unit_Datapath_UA_flag_delay_FFX_4_n1,
         constructing_unit_Datapath_UA_flag_delay_FFX_5_n1,
         constructing_unit_Datapath_UA_flag_delay_FFX_6_n1,
         constructing_unit_Datapath_UA_flag_delay_FFX_7_n1,
         constructing_unit_Datapath_UA_flag_delay_FFX_8_n1,
         constructing_unit_Datapath_UA_flag_delay_FFX_9_n1,
         constructing_unit_Datapath_UA_flag_delay_FFX_10_n1,
         constructing_unit_Datapath_D_h_sq_sample_n1,
         constructing_unit_Datapath_D_v_sq_sample_n4,
         constructing_unit_Datapath_D_v_sq_sample_n3,
         constructing_unit_Datapath_D_v_sq_sample_n2,
         constructing_unit_Datapath_D_v_sq_sample_n1,
         constructing_unit_Datapath_D_adder_add_19_n1,
         constructing_unit_Datapath_D_Cur_tmp_sample_n1,
         constructing_unit_Datapath_D_D_register_n4,
         constructing_unit_Datapath_D_D_register_n3,
         constructing_unit_Datapath_D_D_register_n2,
         constructing_unit_Datapath_D_D_register_n1,
         constructing_unit_Datapath_D_min_register_n92,
         constructing_unit_Datapath_D_min_register_n91,
         constructing_unit_Datapath_D_min_register_n90,
         constructing_unit_Datapath_D_min_register_n89,
         constructing_unit_Datapath_D_min_register_n88,
         constructing_unit_Datapath_D_min_register_n87,
         constructing_unit_Datapath_D_min_register_n86,
         constructing_unit_Datapath_D_min_register_n84,
         constructing_unit_Datapath_D_min_register_n85,
         constructing_unit_Datapath_D_min_register_n83,
         constructing_unit_Datapath_D_min_register_n82,
         constructing_unit_Datapath_D_min_register_n81,
         constructing_unit_Datapath_D_min_register_n80,
         constructing_unit_Datapath_D_min_register_n79,
         constructing_unit_Datapath_D_min_register_n78,
         constructing_unit_Datapath_D_min_register_n77,
         constructing_unit_Datapath_D_min_register_n76,
         constructing_unit_Datapath_D_min_register_n75,
         constructing_unit_Datapath_D_min_register_n74,
         constructing_unit_Datapath_D_min_register_n73,
         constructing_unit_Datapath_D_min_register_n72,
         constructing_unit_Datapath_D_min_register_n71,
         constructing_unit_Datapath_D_min_register_n70,
         constructing_unit_Datapath_D_min_register_n69,
         constructing_unit_Datapath_D_min_register_n68,
         constructing_unit_Datapath_D_min_register_n67,
         constructing_unit_Datapath_D_min_register_n66,
         constructing_unit_Datapath_D_min_register_n65,
         constructing_unit_Datapath_D_min_register_n64,
         constructing_unit_Datapath_D_min_register_n63,
         constructing_unit_Datapath_D_min_register_n62,
         constructing_unit_Datapath_D_min_register_n61,
         constructing_unit_Datapath_D_min_register_n60,
         constructing_unit_Datapath_D_min_register_n59,
         constructing_unit_Datapath_D_min_register_n58,
         constructing_unit_Datapath_D_min_register_n57,
         constructing_unit_Datapath_D_min_register_n56,
         constructing_unit_Datapath_D_min_register_n55,
         constructing_unit_Datapath_D_min_register_n54,
         constructing_unit_Datapath_D_min_register_n53,
         constructing_unit_Datapath_D_min_register_n52,
         constructing_unit_Datapath_D_min_register_n51,
         constructing_unit_Datapath_D_min_register_n50,
         constructing_unit_Datapath_D_min_register_n49,
         constructing_unit_Datapath_D_min_register_n48,
         constructing_unit_Datapath_D_min_register_n47,
         constructing_unit_Datapath_D_min_register_n46,
         constructing_unit_Datapath_D_min_register_n45,
         constructing_unit_Datapath_D_min_register_n44,
         constructing_unit_Datapath_D_min_register_n43,
         constructing_unit_Datapath_D_min_register_n42,
         constructing_unit_Datapath_D_min_register_n41,
         constructing_unit_Datapath_D_min_register_n40,
         constructing_unit_Datapath_D_min_register_n39,
         constructing_unit_Datapath_D_min_register_n38,
         constructing_unit_Datapath_D_min_register_n37,
         constructing_unit_Datapath_D_min_register_n36,
         constructing_unit_Datapath_D_min_register_n35,
         constructing_unit_Datapath_D_min_register_n34,
         constructing_unit_Datapath_D_min_register_n33,
         constructing_unit_Datapath_D_min_register_n32,
         constructing_unit_Datapath_D_min_register_n31,
         constructing_unit_Datapath_D_min_register_n30,
         constructing_unit_Datapath_D_min_register_n29,
         constructing_unit_Datapath_D_min_register_n28,
         constructing_unit_Datapath_D_min_register_n27,
         constructing_unit_Datapath_D_min_register_n26,
         constructing_unit_Datapath_D_min_register_n25,
         constructing_unit_Datapath_D_min_register_n24,
         constructing_unit_Datapath_D_min_register_n23,
         constructing_unit_Datapath_D_min_register_n22,
         constructing_unit_Datapath_D_min_register_n21,
         constructing_unit_Datapath_D_min_register_n20,
         constructing_unit_Datapath_D_min_register_n19,
         constructing_unit_Datapath_D_min_register_n18,
         constructing_unit_Datapath_D_min_register_n17,
         constructing_unit_Datapath_D_min_register_n16,
         constructing_unit_Datapath_D_min_register_n15,
         constructing_unit_Datapath_D_min_register_n14,
         constructing_unit_Datapath_D_min_register_n13,
         constructing_unit_Datapath_D_min_register_n12,
         constructing_unit_Datapath_D_min_register_n11,
         constructing_unit_Datapath_D_min_register_n10,
         constructing_unit_Datapath_D_min_register_n9,
         constructing_unit_Datapath_D_min_register_n8,
         constructing_unit_Datapath_D_min_register_n7,
         constructing_unit_Datapath_D_min_register_n6,
         constructing_unit_Datapath_D_min_register_n5,
         constructing_unit_Datapath_D_min_register_n4,
         constructing_unit_Datapath_D_min_register_n3,
         constructing_unit_Datapath_D_min_register_n2,
         constructing_unit_Datapath_D_min_register_n1,
         constructing_unit_Datapath_final_comp_lt_gt_13_n305,
         constructing_unit_Datapath_final_comp_lt_gt_13_n304,
         constructing_unit_Datapath_final_comp_lt_gt_13_n303,
         constructing_unit_Datapath_final_comp_lt_gt_13_n302,
         constructing_unit_Datapath_final_comp_lt_gt_13_n301,
         constructing_unit_Datapath_final_comp_lt_gt_13_n300,
         constructing_unit_Datapath_final_comp_lt_gt_13_n299,
         constructing_unit_Datapath_final_comp_lt_gt_13_n298,
         constructing_unit_Datapath_final_comp_lt_gt_13_n297,
         constructing_unit_Datapath_final_comp_lt_gt_13_n296,
         constructing_unit_Datapath_final_comp_lt_gt_13_n295,
         constructing_unit_Datapath_final_comp_lt_gt_13_n294,
         constructing_unit_Datapath_final_comp_lt_gt_13_n293,
         constructing_unit_Datapath_final_comp_lt_gt_13_n292,
         constructing_unit_Datapath_final_comp_lt_gt_13_n291,
         constructing_unit_Datapath_final_comp_lt_gt_13_n290,
         constructing_unit_Datapath_final_comp_lt_gt_13_n289,
         constructing_unit_Datapath_final_comp_lt_gt_13_n288,
         constructing_unit_Datapath_final_comp_lt_gt_13_n287,
         constructing_unit_Datapath_final_comp_lt_gt_13_n286,
         constructing_unit_Datapath_final_comp_lt_gt_13_n285,
         constructing_unit_Datapath_final_comp_lt_gt_13_n284,
         constructing_unit_Datapath_final_comp_lt_gt_13_n283,
         constructing_unit_Datapath_final_comp_lt_gt_13_n282,
         constructing_unit_Datapath_final_comp_lt_gt_13_n281,
         constructing_unit_Datapath_final_comp_lt_gt_13_n280,
         constructing_unit_Datapath_final_comp_lt_gt_13_n279,
         constructing_unit_Datapath_final_comp_lt_gt_13_n278,
         constructing_unit_Datapath_final_comp_lt_gt_13_n277,
         constructing_unit_Datapath_final_comp_lt_gt_13_n276,
         constructing_unit_Datapath_final_comp_lt_gt_13_n275,
         constructing_unit_Datapath_final_comp_lt_gt_13_n274,
         constructing_unit_Datapath_final_comp_lt_gt_13_n273,
         constructing_unit_Datapath_final_comp_lt_gt_13_n272,
         constructing_unit_Datapath_final_comp_lt_gt_13_n271,
         constructing_unit_Datapath_final_comp_lt_gt_13_n270,
         constructing_unit_Datapath_final_comp_lt_gt_13_n269,
         constructing_unit_Datapath_final_comp_lt_gt_13_n268,
         constructing_unit_Datapath_final_comp_lt_gt_13_n267,
         constructing_unit_Datapath_final_comp_lt_gt_13_n266,
         constructing_unit_Datapath_final_comp_lt_gt_13_n265,
         constructing_unit_Datapath_final_comp_lt_gt_13_n264,
         constructing_unit_Datapath_final_comp_lt_gt_13_n263,
         constructing_unit_Datapath_final_comp_lt_gt_13_n262,
         constructing_unit_Datapath_final_comp_lt_gt_13_n261,
         constructing_unit_Datapath_final_comp_lt_gt_13_n260,
         constructing_unit_Datapath_final_comp_lt_gt_13_n259,
         constructing_unit_Datapath_final_comp_lt_gt_13_n258,
         constructing_unit_Datapath_final_comp_lt_gt_13_n257,
         constructing_unit_Datapath_final_comp_lt_gt_13_n256,
         constructing_unit_Datapath_final_comp_lt_gt_13_n255,
         constructing_unit_Datapath_final_comp_lt_gt_13_n254,
         constructing_unit_Datapath_final_comp_lt_gt_13_n253,
         constructing_unit_Datapath_final_comp_lt_gt_13_n252,
         constructing_unit_Datapath_final_comp_lt_gt_13_n251,
         constructing_unit_Datapath_final_comp_lt_gt_13_n250,
         constructing_unit_Datapath_final_comp_lt_gt_13_n249,
         constructing_unit_Datapath_final_comp_lt_gt_13_n248,
         constructing_unit_Datapath_final_comp_lt_gt_13_n247,
         constructing_unit_Datapath_final_comp_lt_gt_13_n246,
         constructing_unit_Datapath_final_comp_lt_gt_13_n245,
         constructing_unit_Datapath_final_comp_lt_gt_13_n244,
         constructing_unit_Datapath_final_comp_lt_gt_13_n243,
         constructing_unit_Datapath_final_comp_lt_gt_13_n242,
         constructing_unit_Datapath_final_comp_lt_gt_13_n241,
         constructing_unit_Datapath_final_comp_lt_gt_13_n240,
         constructing_unit_Datapath_final_comp_lt_gt_13_n239,
         constructing_unit_Datapath_final_comp_lt_gt_13_n238,
         constructing_unit_Datapath_final_comp_lt_gt_13_n237,
         constructing_unit_Datapath_final_comp_lt_gt_13_n236,
         constructing_unit_Datapath_final_comp_lt_gt_13_n235,
         constructing_unit_Datapath_final_comp_lt_gt_13_n234,
         constructing_unit_Datapath_final_comp_lt_gt_13_n233,
         constructing_unit_Datapath_final_comp_lt_gt_13_n232,
         constructing_unit_Datapath_final_comp_lt_gt_13_n231,
         constructing_unit_Datapath_final_comp_lt_gt_13_n230,
         constructing_unit_Datapath_final_comp_lt_gt_13_n229,
         constructing_unit_Datapath_final_comp_lt_gt_13_n228,
         constructing_unit_Datapath_final_comp_lt_gt_13_n227,
         constructing_unit_Datapath_final_comp_lt_gt_13_n226,
         constructing_unit_Datapath_final_comp_lt_gt_13_n225,
         constructing_unit_Datapath_final_comp_lt_gt_13_n224,
         constructing_unit_Datapath_final_comp_lt_gt_13_n223,
         constructing_unit_Datapath_final_comp_lt_gt_13_n222,
         constructing_unit_Datapath_final_comp_lt_gt_13_n221,
         constructing_unit_Datapath_final_comp_lt_gt_13_n220,
         constructing_unit_Datapath_final_comp_lt_gt_13_n219,
         constructing_unit_Datapath_final_comp_lt_gt_13_n218,
         constructing_unit_Datapath_final_comp_lt_gt_13_n217,
         constructing_unit_Datapath_final_comp_lt_gt_13_n216,
         constructing_unit_Datapath_final_comp_lt_gt_13_n215,
         constructing_unit_Datapath_final_comp_lt_gt_13_n214,
         constructing_unit_Datapath_final_comp_lt_gt_13_n213,
         constructing_unit_Datapath_final_comp_lt_gt_13_n212,
         constructing_unit_Datapath_final_comp_lt_gt_13_n211,
         constructing_unit_Datapath_final_comp_lt_gt_13_n210,
         constructing_unit_Datapath_final_comp_lt_gt_13_n209,
         constructing_unit_Datapath_final_comp_lt_gt_13_n208,
         constructing_unit_Datapath_final_comp_lt_gt_13_n207,
         constructing_unit_Datapath_final_comp_lt_gt_13_n206,
         constructing_unit_Datapath_final_comp_lt_gt_13_n205,
         constructing_unit_Datapath_final_comp_lt_gt_13_n204,
         constructing_unit_Datapath_final_comp_lt_gt_13_n203,
         constructing_unit_Datapath_final_comp_lt_gt_13_n202,
         constructing_unit_Datapath_final_comp_lt_gt_13_n201,
         constructing_unit_Datapath_final_comp_lt_gt_13_n200,
         constructing_unit_Datapath_comp_out_d_ff_n1,
         constructing_unit_Datapath_COUNT_compEN_n10,
         constructing_unit_Datapath_COUNT_compEN_n8,
         constructing_unit_Datapath_COUNT_compEN_n3,
         constructing_unit_Datapath_COUNT_compEN_n1,
         constructing_unit_Datapath_COUNT_compEN_n9,
         constructing_unit_Datapath_COUNT_compEN_n7,
         constructing_unit_Datapath_COUNT_compEN_n6,
         constructing_unit_Datapath_COUNT_compEN_n5,
         constructing_unit_Datapath_COUNT_compEN_n4,
         constructing_unit_Datapath_COUNT_compEN_n2,
         constructing_unit_Datapath_COUNT_STOPcompEN_n11,
         constructing_unit_Datapath_COUNT_STOPcompEN_n5,
         constructing_unit_Datapath_COUNT_STOPcompEN_n3,
         constructing_unit_Datapath_COUNT_STOPcompEN_n12,
         constructing_unit_Datapath_COUNT_STOPcompEN_n10,
         constructing_unit_Datapath_COUNT_STOPcompEN_n9,
         constructing_unit_Datapath_COUNT_STOPcompEN_n8,
         constructing_unit_Datapath_COUNT_STOPcompEN_n7,
         constructing_unit_Datapath_COUNT_STOPcompEN_n6,
         constructing_unit_Datapath_COUNT_STOPcompEN_n4,
         constructing_unit_Datapath_COUNT_STOPcompEN_n2,
         constructing_unit_Datapath_COUNT_STOPcompEN_n1,
         constructing_unit_Datapath_FaS_registers0_v_1_n33,
         constructing_unit_Datapath_FaS_registers0_v_1_n34,
         constructing_unit_Datapath_FaS_registers0_v_1_n32,
         constructing_unit_Datapath_FaS_registers0_v_1_n31,
         constructing_unit_Datapath_FaS_registers0_v_1_n30,
         constructing_unit_Datapath_FaS_registers0_v_1_n29,
         constructing_unit_Datapath_FaS_registers0_v_1_n28,
         constructing_unit_Datapath_FaS_registers0_v_1_n27,
         constructing_unit_Datapath_FaS_registers0_v_1_n26,
         constructing_unit_Datapath_FaS_registers0_v_1_n25,
         constructing_unit_Datapath_FaS_registers0_v_1_n24,
         constructing_unit_Datapath_FaS_registers0_v_1_n23,
         constructing_unit_Datapath_FaS_registers0_v_1_n22,
         constructing_unit_Datapath_FaS_registers0_v_1_n21,
         constructing_unit_Datapath_FaS_registers0_v_1_n20,
         constructing_unit_Datapath_FaS_registers0_v_1_n19,
         constructing_unit_Datapath_FaS_registers0_v_1_n18,
         constructing_unit_Datapath_FaS_registers0_v_1_n17,
         constructing_unit_Datapath_FaS_registers0_v_1_n16,
         constructing_unit_Datapath_FaS_registers0_v_1_n15,
         constructing_unit_Datapath_FaS_registers0_v_1_n14,
         constructing_unit_Datapath_FaS_registers0_v_1_n13,
         constructing_unit_Datapath_FaS_registers0_v_1_n12,
         constructing_unit_Datapath_FaS_registers0_v_1_n11,
         constructing_unit_Datapath_FaS_registers0_v_1_n10,
         constructing_unit_Datapath_FaS_registers0_v_1_n9,
         constructing_unit_Datapath_FaS_registers0_v_1_n8,
         constructing_unit_Datapath_FaS_registers0_v_1_n7,
         constructing_unit_Datapath_FaS_registers0_v_1_n6,
         constructing_unit_Datapath_FaS_registers0_v_1_n5,
         constructing_unit_Datapath_FaS_registers0_v_1_n4,
         constructing_unit_Datapath_FaS_registers0_v_1_n3,
         constructing_unit_Datapath_FaS_registers0_v_1_n2,
         constructing_unit_Datapath_FaS_registers0_v_1_n1,
         constructing_unit_Datapath_FaS_registers0_v_2_n67,
         constructing_unit_Datapath_FaS_registers0_v_2_n66,
         constructing_unit_Datapath_FaS_registers0_v_2_n65,
         constructing_unit_Datapath_FaS_registers0_v_2_n64,
         constructing_unit_Datapath_FaS_registers0_v_2_n63,
         constructing_unit_Datapath_FaS_registers0_v_2_n62,
         constructing_unit_Datapath_FaS_registers0_v_2_n61,
         constructing_unit_Datapath_FaS_registers0_v_2_n60,
         constructing_unit_Datapath_FaS_registers0_v_2_n59,
         constructing_unit_Datapath_FaS_registers0_v_2_n58,
         constructing_unit_Datapath_FaS_registers0_v_2_n57,
         constructing_unit_Datapath_FaS_registers0_v_2_n56,
         constructing_unit_Datapath_FaS_registers0_v_2_n55,
         constructing_unit_Datapath_FaS_registers0_v_2_n54,
         constructing_unit_Datapath_FaS_registers0_v_2_n53,
         constructing_unit_Datapath_FaS_registers0_v_2_n52,
         constructing_unit_Datapath_FaS_registers0_v_2_n51,
         constructing_unit_Datapath_FaS_registers0_v_2_n50,
         constructing_unit_Datapath_FaS_registers0_v_2_n49,
         constructing_unit_Datapath_FaS_registers0_v_2_n48,
         constructing_unit_Datapath_FaS_registers0_v_2_n47,
         constructing_unit_Datapath_FaS_registers0_v_2_n46,
         constructing_unit_Datapath_FaS_registers0_v_2_n45,
         constructing_unit_Datapath_FaS_registers0_v_2_n44,
         constructing_unit_Datapath_FaS_registers0_v_2_n43,
         constructing_unit_Datapath_FaS_registers0_v_2_n42,
         constructing_unit_Datapath_FaS_registers0_v_2_n41,
         constructing_unit_Datapath_FaS_registers0_v_2_n40,
         constructing_unit_Datapath_FaS_registers0_v_2_n39,
         constructing_unit_Datapath_FaS_registers0_v_2_n38,
         constructing_unit_Datapath_FaS_registers0_v_2_n37,
         constructing_unit_Datapath_FaS_registers0_v_2_n36,
         constructing_unit_Datapath_FaS_registers0_v_2_n35,
         constructing_unit_Datapath_FaS_registers0_v_2_n33,
         constructing_unit_Datapath_FaS_registers1_v_1_n67,
         constructing_unit_Datapath_FaS_registers1_v_1_n66,
         constructing_unit_Datapath_FaS_registers1_v_1_n65,
         constructing_unit_Datapath_FaS_registers1_v_1_n64,
         constructing_unit_Datapath_FaS_registers1_v_1_n63,
         constructing_unit_Datapath_FaS_registers1_v_1_n62,
         constructing_unit_Datapath_FaS_registers1_v_1_n61,
         constructing_unit_Datapath_FaS_registers1_v_1_n60,
         constructing_unit_Datapath_FaS_registers1_v_1_n59,
         constructing_unit_Datapath_FaS_registers1_v_1_n58,
         constructing_unit_Datapath_FaS_registers1_v_1_n57,
         constructing_unit_Datapath_FaS_registers1_v_1_n56,
         constructing_unit_Datapath_FaS_registers1_v_1_n55,
         constructing_unit_Datapath_FaS_registers1_v_1_n54,
         constructing_unit_Datapath_FaS_registers1_v_1_n53,
         constructing_unit_Datapath_FaS_registers1_v_1_n52,
         constructing_unit_Datapath_FaS_registers1_v_1_n51,
         constructing_unit_Datapath_FaS_registers1_v_1_n50,
         constructing_unit_Datapath_FaS_registers1_v_1_n49,
         constructing_unit_Datapath_FaS_registers1_v_1_n48,
         constructing_unit_Datapath_FaS_registers1_v_1_n47,
         constructing_unit_Datapath_FaS_registers1_v_1_n46,
         constructing_unit_Datapath_FaS_registers1_v_1_n45,
         constructing_unit_Datapath_FaS_registers1_v_1_n44,
         constructing_unit_Datapath_FaS_registers1_v_1_n43,
         constructing_unit_Datapath_FaS_registers1_v_1_n42,
         constructing_unit_Datapath_FaS_registers1_v_1_n41,
         constructing_unit_Datapath_FaS_registers1_v_1_n40,
         constructing_unit_Datapath_FaS_registers1_v_1_n39,
         constructing_unit_Datapath_FaS_registers1_v_1_n38,
         constructing_unit_Datapath_FaS_registers1_v_1_n37,
         constructing_unit_Datapath_FaS_registers1_v_1_n36,
         constructing_unit_Datapath_FaS_registers1_v_1_n35,
         constructing_unit_Datapath_FaS_registers1_v_1_n33,
         constructing_unit_Datapath_FaS_registers1_v_2_n67,
         constructing_unit_Datapath_FaS_registers1_v_2_n66,
         constructing_unit_Datapath_FaS_registers1_v_2_n65,
         constructing_unit_Datapath_FaS_registers1_v_2_n64,
         constructing_unit_Datapath_FaS_registers1_v_2_n63,
         constructing_unit_Datapath_FaS_registers1_v_2_n62,
         constructing_unit_Datapath_FaS_registers1_v_2_n61,
         constructing_unit_Datapath_FaS_registers1_v_2_n60,
         constructing_unit_Datapath_FaS_registers1_v_2_n59,
         constructing_unit_Datapath_FaS_registers1_v_2_n58,
         constructing_unit_Datapath_FaS_registers1_v_2_n57,
         constructing_unit_Datapath_FaS_registers1_v_2_n56,
         constructing_unit_Datapath_FaS_registers1_v_2_n55,
         constructing_unit_Datapath_FaS_registers1_v_2_n54,
         constructing_unit_Datapath_FaS_registers1_v_2_n53,
         constructing_unit_Datapath_FaS_registers1_v_2_n52,
         constructing_unit_Datapath_FaS_registers1_v_2_n51,
         constructing_unit_Datapath_FaS_registers1_v_2_n50,
         constructing_unit_Datapath_FaS_registers1_v_2_n49,
         constructing_unit_Datapath_FaS_registers1_v_2_n48,
         constructing_unit_Datapath_FaS_registers1_v_2_n47,
         constructing_unit_Datapath_FaS_registers1_v_2_n46,
         constructing_unit_Datapath_FaS_registers1_v_2_n45,
         constructing_unit_Datapath_FaS_registers1_v_2_n44,
         constructing_unit_Datapath_FaS_registers1_v_2_n43,
         constructing_unit_Datapath_FaS_registers1_v_2_n42,
         constructing_unit_Datapath_FaS_registers1_v_2_n41,
         constructing_unit_Datapath_FaS_registers1_v_2_n40,
         constructing_unit_Datapath_FaS_registers1_v_2_n39,
         constructing_unit_Datapath_FaS_registers1_v_2_n38,
         constructing_unit_Datapath_FaS_registers1_v_2_n37,
         constructing_unit_Datapath_FaS_registers1_v_2_n36,
         constructing_unit_Datapath_FaS_registers1_v_2_n35,
         constructing_unit_Datapath_FaS_registers1_v_2_n33,
         constructing_unit_Datapath_FaS_registers2_v_1_n67,
         constructing_unit_Datapath_FaS_registers2_v_1_n66,
         constructing_unit_Datapath_FaS_registers2_v_1_n65,
         constructing_unit_Datapath_FaS_registers2_v_1_n64,
         constructing_unit_Datapath_FaS_registers2_v_1_n63,
         constructing_unit_Datapath_FaS_registers2_v_1_n62,
         constructing_unit_Datapath_FaS_registers2_v_1_n61,
         constructing_unit_Datapath_FaS_registers2_v_1_n60,
         constructing_unit_Datapath_FaS_registers2_v_1_n59,
         constructing_unit_Datapath_FaS_registers2_v_1_n58,
         constructing_unit_Datapath_FaS_registers2_v_1_n57,
         constructing_unit_Datapath_FaS_registers2_v_1_n56,
         constructing_unit_Datapath_FaS_registers2_v_1_n55,
         constructing_unit_Datapath_FaS_registers2_v_1_n54,
         constructing_unit_Datapath_FaS_registers2_v_1_n53,
         constructing_unit_Datapath_FaS_registers2_v_1_n52,
         constructing_unit_Datapath_FaS_registers2_v_1_n51,
         constructing_unit_Datapath_FaS_registers2_v_1_n50,
         constructing_unit_Datapath_FaS_registers2_v_1_n49,
         constructing_unit_Datapath_FaS_registers2_v_1_n48,
         constructing_unit_Datapath_FaS_registers2_v_1_n47,
         constructing_unit_Datapath_FaS_registers2_v_1_n46,
         constructing_unit_Datapath_FaS_registers2_v_1_n45,
         constructing_unit_Datapath_FaS_registers2_v_1_n44,
         constructing_unit_Datapath_FaS_registers2_v_1_n43,
         constructing_unit_Datapath_FaS_registers2_v_1_n42,
         constructing_unit_Datapath_FaS_registers2_v_1_n41,
         constructing_unit_Datapath_FaS_registers2_v_1_n40,
         constructing_unit_Datapath_FaS_registers2_v_1_n39,
         constructing_unit_Datapath_FaS_registers2_v_1_n38,
         constructing_unit_Datapath_FaS_registers2_v_1_n37,
         constructing_unit_Datapath_FaS_registers2_v_1_n36,
         constructing_unit_Datapath_FaS_registers2_v_1_n35,
         constructing_unit_Datapath_FaS_registers2_v_1_n33,
         constructing_unit_Datapath_FaS_registers2_v_2_n67,
         constructing_unit_Datapath_FaS_registers2_v_2_n66,
         constructing_unit_Datapath_FaS_registers2_v_2_n65,
         constructing_unit_Datapath_FaS_registers2_v_2_n64,
         constructing_unit_Datapath_FaS_registers2_v_2_n63,
         constructing_unit_Datapath_FaS_registers2_v_2_n62,
         constructing_unit_Datapath_FaS_registers2_v_2_n61,
         constructing_unit_Datapath_FaS_registers2_v_2_n60,
         constructing_unit_Datapath_FaS_registers2_v_2_n59,
         constructing_unit_Datapath_FaS_registers2_v_2_n58,
         constructing_unit_Datapath_FaS_registers2_v_2_n57,
         constructing_unit_Datapath_FaS_registers2_v_2_n56,
         constructing_unit_Datapath_FaS_registers2_v_2_n55,
         constructing_unit_Datapath_FaS_registers2_v_2_n54,
         constructing_unit_Datapath_FaS_registers2_v_2_n53,
         constructing_unit_Datapath_FaS_registers2_v_2_n52,
         constructing_unit_Datapath_FaS_registers2_v_2_n51,
         constructing_unit_Datapath_FaS_registers2_v_2_n50,
         constructing_unit_Datapath_FaS_registers2_v_2_n49,
         constructing_unit_Datapath_FaS_registers2_v_2_n48,
         constructing_unit_Datapath_FaS_registers2_v_2_n47,
         constructing_unit_Datapath_FaS_registers2_v_2_n46,
         constructing_unit_Datapath_FaS_registers2_v_2_n45,
         constructing_unit_Datapath_FaS_registers2_v_2_n44,
         constructing_unit_Datapath_FaS_registers2_v_2_n43,
         constructing_unit_Datapath_FaS_registers2_v_2_n42,
         constructing_unit_Datapath_FaS_registers2_v_2_n41,
         constructing_unit_Datapath_FaS_registers2_v_2_n40,
         constructing_unit_Datapath_FaS_registers2_v_2_n39,
         constructing_unit_Datapath_FaS_registers2_v_2_n38,
         constructing_unit_Datapath_FaS_registers2_v_2_n37,
         constructing_unit_Datapath_FaS_registers2_v_2_n36,
         constructing_unit_Datapath_FaS_registers2_v_2_n35,
         constructing_unit_Datapath_FaS_registers2_v_2_n33,
         constructing_unit_Datapath_Middle_registers0_v_3_n67,
         constructing_unit_Datapath_Middle_registers0_v_3_n66,
         constructing_unit_Datapath_Middle_registers0_v_3_n65,
         constructing_unit_Datapath_Middle_registers0_v_3_n64,
         constructing_unit_Datapath_Middle_registers0_v_3_n63,
         constructing_unit_Datapath_Middle_registers0_v_3_n62,
         constructing_unit_Datapath_Middle_registers0_v_3_n61,
         constructing_unit_Datapath_Middle_registers0_v_3_n60,
         constructing_unit_Datapath_Middle_registers0_v_3_n59,
         constructing_unit_Datapath_Middle_registers0_v_3_n58,
         constructing_unit_Datapath_Middle_registers0_v_3_n57,
         constructing_unit_Datapath_Middle_registers0_v_3_n56,
         constructing_unit_Datapath_Middle_registers0_v_3_n55,
         constructing_unit_Datapath_Middle_registers0_v_3_n54,
         constructing_unit_Datapath_Middle_registers0_v_3_n53,
         constructing_unit_Datapath_Middle_registers0_v_3_n52,
         constructing_unit_Datapath_Middle_registers0_v_3_n51,
         constructing_unit_Datapath_Middle_registers0_v_3_n50,
         constructing_unit_Datapath_Middle_registers0_v_3_n49,
         constructing_unit_Datapath_Middle_registers0_v_3_n48,
         constructing_unit_Datapath_Middle_registers0_v_3_n47,
         constructing_unit_Datapath_Middle_registers0_v_3_n46,
         constructing_unit_Datapath_Middle_registers0_v_3_n45,
         constructing_unit_Datapath_Middle_registers0_v_3_n44,
         constructing_unit_Datapath_Middle_registers0_v_3_n43,
         constructing_unit_Datapath_Middle_registers0_v_3_n42,
         constructing_unit_Datapath_Middle_registers0_v_3_n41,
         constructing_unit_Datapath_Middle_registers0_v_3_n40,
         constructing_unit_Datapath_Middle_registers0_v_3_n39,
         constructing_unit_Datapath_Middle_registers0_v_3_n38,
         constructing_unit_Datapath_Middle_registers0_v_3_n37,
         constructing_unit_Datapath_Middle_registers0_v_3_n36,
         constructing_unit_Datapath_Middle_registers0_v_3_n35,
         constructing_unit_Datapath_Middle_registers0_v_3_n33,
         constructing_unit_Datapath_Middle_registers0_v_4_n67,
         constructing_unit_Datapath_Middle_registers0_v_4_n66,
         constructing_unit_Datapath_Middle_registers0_v_4_n65,
         constructing_unit_Datapath_Middle_registers0_v_4_n64,
         constructing_unit_Datapath_Middle_registers0_v_4_n63,
         constructing_unit_Datapath_Middle_registers0_v_4_n62,
         constructing_unit_Datapath_Middle_registers0_v_4_n61,
         constructing_unit_Datapath_Middle_registers0_v_4_n60,
         constructing_unit_Datapath_Middle_registers0_v_4_n59,
         constructing_unit_Datapath_Middle_registers0_v_4_n58,
         constructing_unit_Datapath_Middle_registers0_v_4_n57,
         constructing_unit_Datapath_Middle_registers0_v_4_n56,
         constructing_unit_Datapath_Middle_registers0_v_4_n55,
         constructing_unit_Datapath_Middle_registers0_v_4_n54,
         constructing_unit_Datapath_Middle_registers0_v_4_n53,
         constructing_unit_Datapath_Middle_registers0_v_4_n52,
         constructing_unit_Datapath_Middle_registers0_v_4_n51,
         constructing_unit_Datapath_Middle_registers0_v_4_n50,
         constructing_unit_Datapath_Middle_registers0_v_4_n49,
         constructing_unit_Datapath_Middle_registers0_v_4_n48,
         constructing_unit_Datapath_Middle_registers0_v_4_n47,
         constructing_unit_Datapath_Middle_registers0_v_4_n46,
         constructing_unit_Datapath_Middle_registers0_v_4_n45,
         constructing_unit_Datapath_Middle_registers0_v_4_n44,
         constructing_unit_Datapath_Middle_registers0_v_4_n43,
         constructing_unit_Datapath_Middle_registers0_v_4_n42,
         constructing_unit_Datapath_Middle_registers0_v_4_n41,
         constructing_unit_Datapath_Middle_registers0_v_4_n40,
         constructing_unit_Datapath_Middle_registers0_v_4_n39,
         constructing_unit_Datapath_Middle_registers0_v_4_n38,
         constructing_unit_Datapath_Middle_registers0_v_4_n37,
         constructing_unit_Datapath_Middle_registers0_v_4_n36,
         constructing_unit_Datapath_Middle_registers0_v_4_n35,
         constructing_unit_Datapath_Middle_registers0_v_4_n33,
         constructing_unit_Datapath_Middle_registers0_v_5_n67,
         constructing_unit_Datapath_Middle_registers0_v_5_n66,
         constructing_unit_Datapath_Middle_registers0_v_5_n65,
         constructing_unit_Datapath_Middle_registers0_v_5_n64,
         constructing_unit_Datapath_Middle_registers0_v_5_n63,
         constructing_unit_Datapath_Middle_registers0_v_5_n62,
         constructing_unit_Datapath_Middle_registers0_v_5_n61,
         constructing_unit_Datapath_Middle_registers0_v_5_n60,
         constructing_unit_Datapath_Middle_registers0_v_5_n59,
         constructing_unit_Datapath_Middle_registers0_v_5_n58,
         constructing_unit_Datapath_Middle_registers0_v_5_n57,
         constructing_unit_Datapath_Middle_registers0_v_5_n56,
         constructing_unit_Datapath_Middle_registers0_v_5_n55,
         constructing_unit_Datapath_Middle_registers0_v_5_n54,
         constructing_unit_Datapath_Middle_registers0_v_5_n53,
         constructing_unit_Datapath_Middle_registers0_v_5_n52,
         constructing_unit_Datapath_Middle_registers0_v_5_n51,
         constructing_unit_Datapath_Middle_registers0_v_5_n50,
         constructing_unit_Datapath_Middle_registers0_v_5_n49,
         constructing_unit_Datapath_Middle_registers0_v_5_n48,
         constructing_unit_Datapath_Middle_registers0_v_5_n47,
         constructing_unit_Datapath_Middle_registers0_v_5_n46,
         constructing_unit_Datapath_Middle_registers0_v_5_n45,
         constructing_unit_Datapath_Middle_registers0_v_5_n44,
         constructing_unit_Datapath_Middle_registers0_v_5_n43,
         constructing_unit_Datapath_Middle_registers0_v_5_n42,
         constructing_unit_Datapath_Middle_registers0_v_5_n41,
         constructing_unit_Datapath_Middle_registers0_v_5_n40,
         constructing_unit_Datapath_Middle_registers0_v_5_n39,
         constructing_unit_Datapath_Middle_registers0_v_5_n38,
         constructing_unit_Datapath_Middle_registers0_v_5_n37,
         constructing_unit_Datapath_Middle_registers0_v_5_n36,
         constructing_unit_Datapath_Middle_registers0_v_5_n35,
         constructing_unit_Datapath_Middle_registers0_v_5_n33,
         constructing_unit_Datapath_Middle_registers0_v_6_n67,
         constructing_unit_Datapath_Middle_registers0_v_6_n66,
         constructing_unit_Datapath_Middle_registers0_v_6_n65,
         constructing_unit_Datapath_Middle_registers0_v_6_n64,
         constructing_unit_Datapath_Middle_registers0_v_6_n63,
         constructing_unit_Datapath_Middle_registers0_v_6_n62,
         constructing_unit_Datapath_Middle_registers0_v_6_n61,
         constructing_unit_Datapath_Middle_registers0_v_6_n60,
         constructing_unit_Datapath_Middle_registers0_v_6_n59,
         constructing_unit_Datapath_Middle_registers0_v_6_n58,
         constructing_unit_Datapath_Middle_registers0_v_6_n57,
         constructing_unit_Datapath_Middle_registers0_v_6_n56,
         constructing_unit_Datapath_Middle_registers0_v_6_n55,
         constructing_unit_Datapath_Middle_registers0_v_6_n54,
         constructing_unit_Datapath_Middle_registers0_v_6_n53,
         constructing_unit_Datapath_Middle_registers0_v_6_n52,
         constructing_unit_Datapath_Middle_registers0_v_6_n51,
         constructing_unit_Datapath_Middle_registers0_v_6_n50,
         constructing_unit_Datapath_Middle_registers0_v_6_n49,
         constructing_unit_Datapath_Middle_registers0_v_6_n48,
         constructing_unit_Datapath_Middle_registers0_v_6_n47,
         constructing_unit_Datapath_Middle_registers0_v_6_n46,
         constructing_unit_Datapath_Middle_registers0_v_6_n45,
         constructing_unit_Datapath_Middle_registers0_v_6_n44,
         constructing_unit_Datapath_Middle_registers0_v_6_n43,
         constructing_unit_Datapath_Middle_registers0_v_6_n42,
         constructing_unit_Datapath_Middle_registers0_v_6_n41,
         constructing_unit_Datapath_Middle_registers0_v_6_n40,
         constructing_unit_Datapath_Middle_registers0_v_6_n39,
         constructing_unit_Datapath_Middle_registers0_v_6_n38,
         constructing_unit_Datapath_Middle_registers0_v_6_n37,
         constructing_unit_Datapath_Middle_registers0_v_6_n36,
         constructing_unit_Datapath_Middle_registers0_v_6_n35,
         constructing_unit_Datapath_Middle_registers0_v_6_n33,
         constructing_unit_Datapath_Middle_registers0_v_7_n67,
         constructing_unit_Datapath_Middle_registers0_v_7_n66,
         constructing_unit_Datapath_Middle_registers0_v_7_n65,
         constructing_unit_Datapath_Middle_registers0_v_7_n64,
         constructing_unit_Datapath_Middle_registers0_v_7_n63,
         constructing_unit_Datapath_Middle_registers0_v_7_n62,
         constructing_unit_Datapath_Middle_registers0_v_7_n61,
         constructing_unit_Datapath_Middle_registers0_v_7_n60,
         constructing_unit_Datapath_Middle_registers0_v_7_n59,
         constructing_unit_Datapath_Middle_registers0_v_7_n58,
         constructing_unit_Datapath_Middle_registers0_v_7_n57,
         constructing_unit_Datapath_Middle_registers0_v_7_n56,
         constructing_unit_Datapath_Middle_registers0_v_7_n55,
         constructing_unit_Datapath_Middle_registers0_v_7_n54,
         constructing_unit_Datapath_Middle_registers0_v_7_n53,
         constructing_unit_Datapath_Middle_registers0_v_7_n52,
         constructing_unit_Datapath_Middle_registers0_v_7_n51,
         constructing_unit_Datapath_Middle_registers0_v_7_n50,
         constructing_unit_Datapath_Middle_registers0_v_7_n49,
         constructing_unit_Datapath_Middle_registers0_v_7_n48,
         constructing_unit_Datapath_Middle_registers0_v_7_n47,
         constructing_unit_Datapath_Middle_registers0_v_7_n46,
         constructing_unit_Datapath_Middle_registers0_v_7_n45,
         constructing_unit_Datapath_Middle_registers0_v_7_n44,
         constructing_unit_Datapath_Middle_registers0_v_7_n43,
         constructing_unit_Datapath_Middle_registers0_v_7_n42,
         constructing_unit_Datapath_Middle_registers0_v_7_n41,
         constructing_unit_Datapath_Middle_registers0_v_7_n40,
         constructing_unit_Datapath_Middle_registers0_v_7_n39,
         constructing_unit_Datapath_Middle_registers0_v_7_n38,
         constructing_unit_Datapath_Middle_registers0_v_7_n37,
         constructing_unit_Datapath_Middle_registers0_v_7_n36,
         constructing_unit_Datapath_Middle_registers0_v_7_n35,
         constructing_unit_Datapath_Middle_registers0_v_7_n33,
         constructing_unit_Datapath_Middle_registers0_v_8_n67,
         constructing_unit_Datapath_Middle_registers0_v_8_n66,
         constructing_unit_Datapath_Middle_registers0_v_8_n65,
         constructing_unit_Datapath_Middle_registers0_v_8_n64,
         constructing_unit_Datapath_Middle_registers0_v_8_n63,
         constructing_unit_Datapath_Middle_registers0_v_8_n62,
         constructing_unit_Datapath_Middle_registers0_v_8_n61,
         constructing_unit_Datapath_Middle_registers0_v_8_n60,
         constructing_unit_Datapath_Middle_registers0_v_8_n59,
         constructing_unit_Datapath_Middle_registers0_v_8_n58,
         constructing_unit_Datapath_Middle_registers0_v_8_n57,
         constructing_unit_Datapath_Middle_registers0_v_8_n56,
         constructing_unit_Datapath_Middle_registers0_v_8_n55,
         constructing_unit_Datapath_Middle_registers0_v_8_n54,
         constructing_unit_Datapath_Middle_registers0_v_8_n53,
         constructing_unit_Datapath_Middle_registers0_v_8_n52,
         constructing_unit_Datapath_Middle_registers0_v_8_n51,
         constructing_unit_Datapath_Middle_registers0_v_8_n50,
         constructing_unit_Datapath_Middle_registers0_v_8_n49,
         constructing_unit_Datapath_Middle_registers0_v_8_n48,
         constructing_unit_Datapath_Middle_registers0_v_8_n47,
         constructing_unit_Datapath_Middle_registers0_v_8_n46,
         constructing_unit_Datapath_Middle_registers0_v_8_n45,
         constructing_unit_Datapath_Middle_registers0_v_8_n44,
         constructing_unit_Datapath_Middle_registers0_v_8_n43,
         constructing_unit_Datapath_Middle_registers0_v_8_n42,
         constructing_unit_Datapath_Middle_registers0_v_8_n41,
         constructing_unit_Datapath_Middle_registers0_v_8_n40,
         constructing_unit_Datapath_Middle_registers0_v_8_n39,
         constructing_unit_Datapath_Middle_registers0_v_8_n38,
         constructing_unit_Datapath_Middle_registers0_v_8_n37,
         constructing_unit_Datapath_Middle_registers0_v_8_n36,
         constructing_unit_Datapath_Middle_registers0_v_8_n35,
         constructing_unit_Datapath_Middle_registers0_v_8_n33,
         constructing_unit_Datapath_Middle_registers0_v_9_n67,
         constructing_unit_Datapath_Middle_registers0_v_9_n66,
         constructing_unit_Datapath_Middle_registers0_v_9_n65,
         constructing_unit_Datapath_Middle_registers0_v_9_n64,
         constructing_unit_Datapath_Middle_registers0_v_9_n63,
         constructing_unit_Datapath_Middle_registers0_v_9_n62,
         constructing_unit_Datapath_Middle_registers0_v_9_n61,
         constructing_unit_Datapath_Middle_registers0_v_9_n60,
         constructing_unit_Datapath_Middle_registers0_v_9_n59,
         constructing_unit_Datapath_Middle_registers0_v_9_n58,
         constructing_unit_Datapath_Middle_registers0_v_9_n57,
         constructing_unit_Datapath_Middle_registers0_v_9_n56,
         constructing_unit_Datapath_Middle_registers0_v_9_n55,
         constructing_unit_Datapath_Middle_registers0_v_9_n54,
         constructing_unit_Datapath_Middle_registers0_v_9_n53,
         constructing_unit_Datapath_Middle_registers0_v_9_n52,
         constructing_unit_Datapath_Middle_registers0_v_9_n51,
         constructing_unit_Datapath_Middle_registers0_v_9_n50,
         constructing_unit_Datapath_Middle_registers0_v_9_n49,
         constructing_unit_Datapath_Middle_registers0_v_9_n48,
         constructing_unit_Datapath_Middle_registers0_v_9_n47,
         constructing_unit_Datapath_Middle_registers0_v_9_n46,
         constructing_unit_Datapath_Middle_registers0_v_9_n45,
         constructing_unit_Datapath_Middle_registers0_v_9_n44,
         constructing_unit_Datapath_Middle_registers0_v_9_n43,
         constructing_unit_Datapath_Middle_registers0_v_9_n42,
         constructing_unit_Datapath_Middle_registers0_v_9_n41,
         constructing_unit_Datapath_Middle_registers0_v_9_n40,
         constructing_unit_Datapath_Middle_registers0_v_9_n39,
         constructing_unit_Datapath_Middle_registers0_v_9_n38,
         constructing_unit_Datapath_Middle_registers0_v_9_n37,
         constructing_unit_Datapath_Middle_registers0_v_9_n36,
         constructing_unit_Datapath_Middle_registers0_v_9_n35,
         constructing_unit_Datapath_Middle_registers0_v_9_n33,
         constructing_unit_Datapath_Middle_registers0_v_10_n67,
         constructing_unit_Datapath_Middle_registers0_v_10_n66,
         constructing_unit_Datapath_Middle_registers0_v_10_n65,
         constructing_unit_Datapath_Middle_registers0_v_10_n64,
         constructing_unit_Datapath_Middle_registers0_v_10_n63,
         constructing_unit_Datapath_Middle_registers0_v_10_n62,
         constructing_unit_Datapath_Middle_registers0_v_10_n61,
         constructing_unit_Datapath_Middle_registers0_v_10_n60,
         constructing_unit_Datapath_Middle_registers0_v_10_n59,
         constructing_unit_Datapath_Middle_registers0_v_10_n58,
         constructing_unit_Datapath_Middle_registers0_v_10_n57,
         constructing_unit_Datapath_Middle_registers0_v_10_n56,
         constructing_unit_Datapath_Middle_registers0_v_10_n55,
         constructing_unit_Datapath_Middle_registers0_v_10_n54,
         constructing_unit_Datapath_Middle_registers0_v_10_n53,
         constructing_unit_Datapath_Middle_registers0_v_10_n52,
         constructing_unit_Datapath_Middle_registers0_v_10_n51,
         constructing_unit_Datapath_Middle_registers0_v_10_n50,
         constructing_unit_Datapath_Middle_registers0_v_10_n49,
         constructing_unit_Datapath_Middle_registers0_v_10_n48,
         constructing_unit_Datapath_Middle_registers0_v_10_n47,
         constructing_unit_Datapath_Middle_registers0_v_10_n46,
         constructing_unit_Datapath_Middle_registers0_v_10_n45,
         constructing_unit_Datapath_Middle_registers0_v_10_n44,
         constructing_unit_Datapath_Middle_registers0_v_10_n43,
         constructing_unit_Datapath_Middle_registers0_v_10_n42,
         constructing_unit_Datapath_Middle_registers0_v_10_n41,
         constructing_unit_Datapath_Middle_registers0_v_10_n40,
         constructing_unit_Datapath_Middle_registers0_v_10_n39,
         constructing_unit_Datapath_Middle_registers0_v_10_n38,
         constructing_unit_Datapath_Middle_registers0_v_10_n37,
         constructing_unit_Datapath_Middle_registers0_v_10_n36,
         constructing_unit_Datapath_Middle_registers0_v_10_n35,
         constructing_unit_Datapath_Middle_registers0_v_10_n33,
         constructing_unit_Datapath_Middle_registers0_v_11_n67,
         constructing_unit_Datapath_Middle_registers0_v_11_n66,
         constructing_unit_Datapath_Middle_registers0_v_11_n65,
         constructing_unit_Datapath_Middle_registers0_v_11_n64,
         constructing_unit_Datapath_Middle_registers0_v_11_n63,
         constructing_unit_Datapath_Middle_registers0_v_11_n62,
         constructing_unit_Datapath_Middle_registers0_v_11_n61,
         constructing_unit_Datapath_Middle_registers0_v_11_n60,
         constructing_unit_Datapath_Middle_registers0_v_11_n59,
         constructing_unit_Datapath_Middle_registers0_v_11_n58,
         constructing_unit_Datapath_Middle_registers0_v_11_n57,
         constructing_unit_Datapath_Middle_registers0_v_11_n56,
         constructing_unit_Datapath_Middle_registers0_v_11_n55,
         constructing_unit_Datapath_Middle_registers0_v_11_n54,
         constructing_unit_Datapath_Middle_registers0_v_11_n53,
         constructing_unit_Datapath_Middle_registers0_v_11_n52,
         constructing_unit_Datapath_Middle_registers0_v_11_n51,
         constructing_unit_Datapath_Middle_registers0_v_11_n50,
         constructing_unit_Datapath_Middle_registers0_v_11_n49,
         constructing_unit_Datapath_Middle_registers0_v_11_n48,
         constructing_unit_Datapath_Middle_registers0_v_11_n47,
         constructing_unit_Datapath_Middle_registers0_v_11_n46,
         constructing_unit_Datapath_Middle_registers0_v_11_n45,
         constructing_unit_Datapath_Middle_registers0_v_11_n44,
         constructing_unit_Datapath_Middle_registers0_v_11_n43,
         constructing_unit_Datapath_Middle_registers0_v_11_n42,
         constructing_unit_Datapath_Middle_registers0_v_11_n41,
         constructing_unit_Datapath_Middle_registers0_v_11_n40,
         constructing_unit_Datapath_Middle_registers0_v_11_n39,
         constructing_unit_Datapath_Middle_registers0_v_11_n38,
         constructing_unit_Datapath_Middle_registers0_v_11_n37,
         constructing_unit_Datapath_Middle_registers0_v_11_n36,
         constructing_unit_Datapath_Middle_registers0_v_11_n35,
         constructing_unit_Datapath_Middle_registers0_v_11_n33,
         constructing_unit_Datapath_Middle_registers0_v_12_n67,
         constructing_unit_Datapath_Middle_registers0_v_12_n66,
         constructing_unit_Datapath_Middle_registers0_v_12_n65,
         constructing_unit_Datapath_Middle_registers0_v_12_n64,
         constructing_unit_Datapath_Middle_registers0_v_12_n63,
         constructing_unit_Datapath_Middle_registers0_v_12_n62,
         constructing_unit_Datapath_Middle_registers0_v_12_n61,
         constructing_unit_Datapath_Middle_registers0_v_12_n60,
         constructing_unit_Datapath_Middle_registers0_v_12_n59,
         constructing_unit_Datapath_Middle_registers0_v_12_n58,
         constructing_unit_Datapath_Middle_registers0_v_12_n57,
         constructing_unit_Datapath_Middle_registers0_v_12_n56,
         constructing_unit_Datapath_Middle_registers0_v_12_n55,
         constructing_unit_Datapath_Middle_registers0_v_12_n54,
         constructing_unit_Datapath_Middle_registers0_v_12_n53,
         constructing_unit_Datapath_Middle_registers0_v_12_n52,
         constructing_unit_Datapath_Middle_registers0_v_12_n51,
         constructing_unit_Datapath_Middle_registers0_v_12_n50,
         constructing_unit_Datapath_Middle_registers0_v_12_n49,
         constructing_unit_Datapath_Middle_registers0_v_12_n48,
         constructing_unit_Datapath_Middle_registers0_v_12_n47,
         constructing_unit_Datapath_Middle_registers0_v_12_n46,
         constructing_unit_Datapath_Middle_registers0_v_12_n45,
         constructing_unit_Datapath_Middle_registers0_v_12_n44,
         constructing_unit_Datapath_Middle_registers0_v_12_n43,
         constructing_unit_Datapath_Middle_registers0_v_12_n42,
         constructing_unit_Datapath_Middle_registers0_v_12_n41,
         constructing_unit_Datapath_Middle_registers0_v_12_n40,
         constructing_unit_Datapath_Middle_registers0_v_12_n39,
         constructing_unit_Datapath_Middle_registers0_v_12_n38,
         constructing_unit_Datapath_Middle_registers0_v_12_n37,
         constructing_unit_Datapath_Middle_registers0_v_12_n36,
         constructing_unit_Datapath_Middle_registers0_v_12_n35,
         constructing_unit_Datapath_Middle_registers0_v_12_n33,
         constructing_unit_Datapath_Middle_registers0_v_13_n67,
         constructing_unit_Datapath_Middle_registers0_v_13_n66,
         constructing_unit_Datapath_Middle_registers0_v_13_n65,
         constructing_unit_Datapath_Middle_registers0_v_13_n64,
         constructing_unit_Datapath_Middle_registers0_v_13_n63,
         constructing_unit_Datapath_Middle_registers0_v_13_n62,
         constructing_unit_Datapath_Middle_registers0_v_13_n61,
         constructing_unit_Datapath_Middle_registers0_v_13_n60,
         constructing_unit_Datapath_Middle_registers0_v_13_n59,
         constructing_unit_Datapath_Middle_registers0_v_13_n58,
         constructing_unit_Datapath_Middle_registers0_v_13_n57,
         constructing_unit_Datapath_Middle_registers0_v_13_n56,
         constructing_unit_Datapath_Middle_registers0_v_13_n55,
         constructing_unit_Datapath_Middle_registers0_v_13_n54,
         constructing_unit_Datapath_Middle_registers0_v_13_n53,
         constructing_unit_Datapath_Middle_registers0_v_13_n52,
         constructing_unit_Datapath_Middle_registers0_v_13_n51,
         constructing_unit_Datapath_Middle_registers0_v_13_n50,
         constructing_unit_Datapath_Middle_registers0_v_13_n49,
         constructing_unit_Datapath_Middle_registers0_v_13_n48,
         constructing_unit_Datapath_Middle_registers0_v_13_n47,
         constructing_unit_Datapath_Middle_registers0_v_13_n46,
         constructing_unit_Datapath_Middle_registers0_v_13_n45,
         constructing_unit_Datapath_Middle_registers0_v_13_n44,
         constructing_unit_Datapath_Middle_registers0_v_13_n43,
         constructing_unit_Datapath_Middle_registers0_v_13_n42,
         constructing_unit_Datapath_Middle_registers0_v_13_n41,
         constructing_unit_Datapath_Middle_registers0_v_13_n40,
         constructing_unit_Datapath_Middle_registers0_v_13_n39,
         constructing_unit_Datapath_Middle_registers0_v_13_n38,
         constructing_unit_Datapath_Middle_registers0_v_13_n37,
         constructing_unit_Datapath_Middle_registers0_v_13_n36,
         constructing_unit_Datapath_Middle_registers0_v_13_n35,
         constructing_unit_Datapath_Middle_registers0_v_13_n33,
         constructing_unit_Datapath_Middle_registers1_v_3_n67,
         constructing_unit_Datapath_Middle_registers1_v_3_n66,
         constructing_unit_Datapath_Middle_registers1_v_3_n65,
         constructing_unit_Datapath_Middle_registers1_v_3_n64,
         constructing_unit_Datapath_Middle_registers1_v_3_n63,
         constructing_unit_Datapath_Middle_registers1_v_3_n62,
         constructing_unit_Datapath_Middle_registers1_v_3_n61,
         constructing_unit_Datapath_Middle_registers1_v_3_n60,
         constructing_unit_Datapath_Middle_registers1_v_3_n59,
         constructing_unit_Datapath_Middle_registers1_v_3_n58,
         constructing_unit_Datapath_Middle_registers1_v_3_n57,
         constructing_unit_Datapath_Middle_registers1_v_3_n56,
         constructing_unit_Datapath_Middle_registers1_v_3_n55,
         constructing_unit_Datapath_Middle_registers1_v_3_n54,
         constructing_unit_Datapath_Middle_registers1_v_3_n53,
         constructing_unit_Datapath_Middle_registers1_v_3_n52,
         constructing_unit_Datapath_Middle_registers1_v_3_n51,
         constructing_unit_Datapath_Middle_registers1_v_3_n50,
         constructing_unit_Datapath_Middle_registers1_v_3_n49,
         constructing_unit_Datapath_Middle_registers1_v_3_n48,
         constructing_unit_Datapath_Middle_registers1_v_3_n47,
         constructing_unit_Datapath_Middle_registers1_v_3_n46,
         constructing_unit_Datapath_Middle_registers1_v_3_n45,
         constructing_unit_Datapath_Middle_registers1_v_3_n44,
         constructing_unit_Datapath_Middle_registers1_v_3_n43,
         constructing_unit_Datapath_Middle_registers1_v_3_n42,
         constructing_unit_Datapath_Middle_registers1_v_3_n41,
         constructing_unit_Datapath_Middle_registers1_v_3_n40,
         constructing_unit_Datapath_Middle_registers1_v_3_n39,
         constructing_unit_Datapath_Middle_registers1_v_3_n38,
         constructing_unit_Datapath_Middle_registers1_v_3_n37,
         constructing_unit_Datapath_Middle_registers1_v_3_n36,
         constructing_unit_Datapath_Middle_registers1_v_3_n35,
         constructing_unit_Datapath_Middle_registers1_v_3_n33,
         constructing_unit_Datapath_Middle_registers1_v_4_n67,
         constructing_unit_Datapath_Middle_registers1_v_4_n66,
         constructing_unit_Datapath_Middle_registers1_v_4_n65,
         constructing_unit_Datapath_Middle_registers1_v_4_n64,
         constructing_unit_Datapath_Middle_registers1_v_4_n63,
         constructing_unit_Datapath_Middle_registers1_v_4_n62,
         constructing_unit_Datapath_Middle_registers1_v_4_n61,
         constructing_unit_Datapath_Middle_registers1_v_4_n60,
         constructing_unit_Datapath_Middle_registers1_v_4_n59,
         constructing_unit_Datapath_Middle_registers1_v_4_n58,
         constructing_unit_Datapath_Middle_registers1_v_4_n57,
         constructing_unit_Datapath_Middle_registers1_v_4_n56,
         constructing_unit_Datapath_Middle_registers1_v_4_n55,
         constructing_unit_Datapath_Middle_registers1_v_4_n54,
         constructing_unit_Datapath_Middle_registers1_v_4_n53,
         constructing_unit_Datapath_Middle_registers1_v_4_n52,
         constructing_unit_Datapath_Middle_registers1_v_4_n51,
         constructing_unit_Datapath_Middle_registers1_v_4_n50,
         constructing_unit_Datapath_Middle_registers1_v_4_n49,
         constructing_unit_Datapath_Middle_registers1_v_4_n48,
         constructing_unit_Datapath_Middle_registers1_v_4_n47,
         constructing_unit_Datapath_Middle_registers1_v_4_n46,
         constructing_unit_Datapath_Middle_registers1_v_4_n45,
         constructing_unit_Datapath_Middle_registers1_v_4_n44,
         constructing_unit_Datapath_Middle_registers1_v_4_n43,
         constructing_unit_Datapath_Middle_registers1_v_4_n42,
         constructing_unit_Datapath_Middle_registers1_v_4_n41,
         constructing_unit_Datapath_Middle_registers1_v_4_n40,
         constructing_unit_Datapath_Middle_registers1_v_4_n39,
         constructing_unit_Datapath_Middle_registers1_v_4_n38,
         constructing_unit_Datapath_Middle_registers1_v_4_n37,
         constructing_unit_Datapath_Middle_registers1_v_4_n36,
         constructing_unit_Datapath_Middle_registers1_v_4_n35,
         constructing_unit_Datapath_Middle_registers1_v_4_n33,
         constructing_unit_Datapath_Middle_registers1_v_5_n67,
         constructing_unit_Datapath_Middle_registers1_v_5_n66,
         constructing_unit_Datapath_Middle_registers1_v_5_n65,
         constructing_unit_Datapath_Middle_registers1_v_5_n64,
         constructing_unit_Datapath_Middle_registers1_v_5_n63,
         constructing_unit_Datapath_Middle_registers1_v_5_n62,
         constructing_unit_Datapath_Middle_registers1_v_5_n61,
         constructing_unit_Datapath_Middle_registers1_v_5_n60,
         constructing_unit_Datapath_Middle_registers1_v_5_n59,
         constructing_unit_Datapath_Middle_registers1_v_5_n58,
         constructing_unit_Datapath_Middle_registers1_v_5_n57,
         constructing_unit_Datapath_Middle_registers1_v_5_n56,
         constructing_unit_Datapath_Middle_registers1_v_5_n55,
         constructing_unit_Datapath_Middle_registers1_v_5_n54,
         constructing_unit_Datapath_Middle_registers1_v_5_n53,
         constructing_unit_Datapath_Middle_registers1_v_5_n52,
         constructing_unit_Datapath_Middle_registers1_v_5_n51,
         constructing_unit_Datapath_Middle_registers1_v_5_n50,
         constructing_unit_Datapath_Middle_registers1_v_5_n49,
         constructing_unit_Datapath_Middle_registers1_v_5_n48,
         constructing_unit_Datapath_Middle_registers1_v_5_n47,
         constructing_unit_Datapath_Middle_registers1_v_5_n46,
         constructing_unit_Datapath_Middle_registers1_v_5_n45,
         constructing_unit_Datapath_Middle_registers1_v_5_n44,
         constructing_unit_Datapath_Middle_registers1_v_5_n43,
         constructing_unit_Datapath_Middle_registers1_v_5_n42,
         constructing_unit_Datapath_Middle_registers1_v_5_n41,
         constructing_unit_Datapath_Middle_registers1_v_5_n40,
         constructing_unit_Datapath_Middle_registers1_v_5_n39,
         constructing_unit_Datapath_Middle_registers1_v_5_n38,
         constructing_unit_Datapath_Middle_registers1_v_5_n37,
         constructing_unit_Datapath_Middle_registers1_v_5_n36,
         constructing_unit_Datapath_Middle_registers1_v_5_n35,
         constructing_unit_Datapath_Middle_registers1_v_5_n33,
         constructing_unit_Datapath_Middle_registers1_v_6_n67,
         constructing_unit_Datapath_Middle_registers1_v_6_n66,
         constructing_unit_Datapath_Middle_registers1_v_6_n65,
         constructing_unit_Datapath_Middle_registers1_v_6_n64,
         constructing_unit_Datapath_Middle_registers1_v_6_n63,
         constructing_unit_Datapath_Middle_registers1_v_6_n62,
         constructing_unit_Datapath_Middle_registers1_v_6_n61,
         constructing_unit_Datapath_Middle_registers1_v_6_n60,
         constructing_unit_Datapath_Middle_registers1_v_6_n59,
         constructing_unit_Datapath_Middle_registers1_v_6_n58,
         constructing_unit_Datapath_Middle_registers1_v_6_n57,
         constructing_unit_Datapath_Middle_registers1_v_6_n56,
         constructing_unit_Datapath_Middle_registers1_v_6_n55,
         constructing_unit_Datapath_Middle_registers1_v_6_n54,
         constructing_unit_Datapath_Middle_registers1_v_6_n53,
         constructing_unit_Datapath_Middle_registers1_v_6_n52,
         constructing_unit_Datapath_Middle_registers1_v_6_n51,
         constructing_unit_Datapath_Middle_registers1_v_6_n50,
         constructing_unit_Datapath_Middle_registers1_v_6_n49,
         constructing_unit_Datapath_Middle_registers1_v_6_n48,
         constructing_unit_Datapath_Middle_registers1_v_6_n47,
         constructing_unit_Datapath_Middle_registers1_v_6_n46,
         constructing_unit_Datapath_Middle_registers1_v_6_n45,
         constructing_unit_Datapath_Middle_registers1_v_6_n44,
         constructing_unit_Datapath_Middle_registers1_v_6_n43,
         constructing_unit_Datapath_Middle_registers1_v_6_n42,
         constructing_unit_Datapath_Middle_registers1_v_6_n41,
         constructing_unit_Datapath_Middle_registers1_v_6_n40,
         constructing_unit_Datapath_Middle_registers1_v_6_n39,
         constructing_unit_Datapath_Middle_registers1_v_6_n38,
         constructing_unit_Datapath_Middle_registers1_v_6_n37,
         constructing_unit_Datapath_Middle_registers1_v_6_n36,
         constructing_unit_Datapath_Middle_registers1_v_6_n35,
         constructing_unit_Datapath_Middle_registers1_v_6_n33,
         constructing_unit_Datapath_Middle_registers1_v_7_n67,
         constructing_unit_Datapath_Middle_registers1_v_7_n66,
         constructing_unit_Datapath_Middle_registers1_v_7_n65,
         constructing_unit_Datapath_Middle_registers1_v_7_n64,
         constructing_unit_Datapath_Middle_registers1_v_7_n63,
         constructing_unit_Datapath_Middle_registers1_v_7_n62,
         constructing_unit_Datapath_Middle_registers1_v_7_n61,
         constructing_unit_Datapath_Middle_registers1_v_7_n60,
         constructing_unit_Datapath_Middle_registers1_v_7_n59,
         constructing_unit_Datapath_Middle_registers1_v_7_n58,
         constructing_unit_Datapath_Middle_registers1_v_7_n57,
         constructing_unit_Datapath_Middle_registers1_v_7_n56,
         constructing_unit_Datapath_Middle_registers1_v_7_n55,
         constructing_unit_Datapath_Middle_registers1_v_7_n54,
         constructing_unit_Datapath_Middle_registers1_v_7_n53,
         constructing_unit_Datapath_Middle_registers1_v_7_n52,
         constructing_unit_Datapath_Middle_registers1_v_7_n51,
         constructing_unit_Datapath_Middle_registers1_v_7_n50,
         constructing_unit_Datapath_Middle_registers1_v_7_n49,
         constructing_unit_Datapath_Middle_registers1_v_7_n48,
         constructing_unit_Datapath_Middle_registers1_v_7_n47,
         constructing_unit_Datapath_Middle_registers1_v_7_n46,
         constructing_unit_Datapath_Middle_registers1_v_7_n45,
         constructing_unit_Datapath_Middle_registers1_v_7_n44,
         constructing_unit_Datapath_Middle_registers1_v_7_n43,
         constructing_unit_Datapath_Middle_registers1_v_7_n42,
         constructing_unit_Datapath_Middle_registers1_v_7_n41,
         constructing_unit_Datapath_Middle_registers1_v_7_n40,
         constructing_unit_Datapath_Middle_registers1_v_7_n39,
         constructing_unit_Datapath_Middle_registers1_v_7_n38,
         constructing_unit_Datapath_Middle_registers1_v_7_n37,
         constructing_unit_Datapath_Middle_registers1_v_7_n36,
         constructing_unit_Datapath_Middle_registers1_v_7_n35,
         constructing_unit_Datapath_Middle_registers1_v_7_n33,
         constructing_unit_Datapath_Middle_registers1_v_8_n67,
         constructing_unit_Datapath_Middle_registers1_v_8_n66,
         constructing_unit_Datapath_Middle_registers1_v_8_n65,
         constructing_unit_Datapath_Middle_registers1_v_8_n64,
         constructing_unit_Datapath_Middle_registers1_v_8_n63,
         constructing_unit_Datapath_Middle_registers1_v_8_n62,
         constructing_unit_Datapath_Middle_registers1_v_8_n61,
         constructing_unit_Datapath_Middle_registers1_v_8_n60,
         constructing_unit_Datapath_Middle_registers1_v_8_n59,
         constructing_unit_Datapath_Middle_registers1_v_8_n58,
         constructing_unit_Datapath_Middle_registers1_v_8_n57,
         constructing_unit_Datapath_Middle_registers1_v_8_n56,
         constructing_unit_Datapath_Middle_registers1_v_8_n55,
         constructing_unit_Datapath_Middle_registers1_v_8_n54,
         constructing_unit_Datapath_Middle_registers1_v_8_n53,
         constructing_unit_Datapath_Middle_registers1_v_8_n52,
         constructing_unit_Datapath_Middle_registers1_v_8_n51,
         constructing_unit_Datapath_Middle_registers1_v_8_n50,
         constructing_unit_Datapath_Middle_registers1_v_8_n49,
         constructing_unit_Datapath_Middle_registers1_v_8_n48,
         constructing_unit_Datapath_Middle_registers1_v_8_n47,
         constructing_unit_Datapath_Middle_registers1_v_8_n46,
         constructing_unit_Datapath_Middle_registers1_v_8_n45,
         constructing_unit_Datapath_Middle_registers1_v_8_n44,
         constructing_unit_Datapath_Middle_registers1_v_8_n43,
         constructing_unit_Datapath_Middle_registers1_v_8_n42,
         constructing_unit_Datapath_Middle_registers1_v_8_n41,
         constructing_unit_Datapath_Middle_registers1_v_8_n40,
         constructing_unit_Datapath_Middle_registers1_v_8_n39,
         constructing_unit_Datapath_Middle_registers1_v_8_n38,
         constructing_unit_Datapath_Middle_registers1_v_8_n37,
         constructing_unit_Datapath_Middle_registers1_v_8_n36,
         constructing_unit_Datapath_Middle_registers1_v_8_n35,
         constructing_unit_Datapath_Middle_registers1_v_8_n33,
         constructing_unit_Datapath_Middle_registers1_v_9_n67,
         constructing_unit_Datapath_Middle_registers1_v_9_n66,
         constructing_unit_Datapath_Middle_registers1_v_9_n65,
         constructing_unit_Datapath_Middle_registers1_v_9_n64,
         constructing_unit_Datapath_Middle_registers1_v_9_n63,
         constructing_unit_Datapath_Middle_registers1_v_9_n62,
         constructing_unit_Datapath_Middle_registers1_v_9_n61,
         constructing_unit_Datapath_Middle_registers1_v_9_n60,
         constructing_unit_Datapath_Middle_registers1_v_9_n59,
         constructing_unit_Datapath_Middle_registers1_v_9_n58,
         constructing_unit_Datapath_Middle_registers1_v_9_n57,
         constructing_unit_Datapath_Middle_registers1_v_9_n56,
         constructing_unit_Datapath_Middle_registers1_v_9_n55,
         constructing_unit_Datapath_Middle_registers1_v_9_n54,
         constructing_unit_Datapath_Middle_registers1_v_9_n53,
         constructing_unit_Datapath_Middle_registers1_v_9_n52,
         constructing_unit_Datapath_Middle_registers1_v_9_n51,
         constructing_unit_Datapath_Middle_registers1_v_9_n50,
         constructing_unit_Datapath_Middle_registers1_v_9_n49,
         constructing_unit_Datapath_Middle_registers1_v_9_n48,
         constructing_unit_Datapath_Middle_registers1_v_9_n47,
         constructing_unit_Datapath_Middle_registers1_v_9_n46,
         constructing_unit_Datapath_Middle_registers1_v_9_n45,
         constructing_unit_Datapath_Middle_registers1_v_9_n44,
         constructing_unit_Datapath_Middle_registers1_v_9_n43,
         constructing_unit_Datapath_Middle_registers1_v_9_n42,
         constructing_unit_Datapath_Middle_registers1_v_9_n41,
         constructing_unit_Datapath_Middle_registers1_v_9_n40,
         constructing_unit_Datapath_Middle_registers1_v_9_n39,
         constructing_unit_Datapath_Middle_registers1_v_9_n38,
         constructing_unit_Datapath_Middle_registers1_v_9_n37,
         constructing_unit_Datapath_Middle_registers1_v_9_n36,
         constructing_unit_Datapath_Middle_registers1_v_9_n35,
         constructing_unit_Datapath_Middle_registers1_v_9_n33,
         constructing_unit_Datapath_Middle_registers1_v_10_n67,
         constructing_unit_Datapath_Middle_registers1_v_10_n66,
         constructing_unit_Datapath_Middle_registers1_v_10_n65,
         constructing_unit_Datapath_Middle_registers1_v_10_n64,
         constructing_unit_Datapath_Middle_registers1_v_10_n63,
         constructing_unit_Datapath_Middle_registers1_v_10_n62,
         constructing_unit_Datapath_Middle_registers1_v_10_n61,
         constructing_unit_Datapath_Middle_registers1_v_10_n60,
         constructing_unit_Datapath_Middle_registers1_v_10_n59,
         constructing_unit_Datapath_Middle_registers1_v_10_n58,
         constructing_unit_Datapath_Middle_registers1_v_10_n57,
         constructing_unit_Datapath_Middle_registers1_v_10_n56,
         constructing_unit_Datapath_Middle_registers1_v_10_n55,
         constructing_unit_Datapath_Middle_registers1_v_10_n54,
         constructing_unit_Datapath_Middle_registers1_v_10_n53,
         constructing_unit_Datapath_Middle_registers1_v_10_n52,
         constructing_unit_Datapath_Middle_registers1_v_10_n51,
         constructing_unit_Datapath_Middle_registers1_v_10_n50,
         constructing_unit_Datapath_Middle_registers1_v_10_n49,
         constructing_unit_Datapath_Middle_registers1_v_10_n48,
         constructing_unit_Datapath_Middle_registers1_v_10_n47,
         constructing_unit_Datapath_Middle_registers1_v_10_n46,
         constructing_unit_Datapath_Middle_registers1_v_10_n45,
         constructing_unit_Datapath_Middle_registers1_v_10_n44,
         constructing_unit_Datapath_Middle_registers1_v_10_n43,
         constructing_unit_Datapath_Middle_registers1_v_10_n42,
         constructing_unit_Datapath_Middle_registers1_v_10_n41,
         constructing_unit_Datapath_Middle_registers1_v_10_n40,
         constructing_unit_Datapath_Middle_registers1_v_10_n39,
         constructing_unit_Datapath_Middle_registers1_v_10_n38,
         constructing_unit_Datapath_Middle_registers1_v_10_n37,
         constructing_unit_Datapath_Middle_registers1_v_10_n36,
         constructing_unit_Datapath_Middle_registers1_v_10_n35,
         constructing_unit_Datapath_Middle_registers1_v_10_n33,
         constructing_unit_Datapath_Middle_registers1_v_11_n67,
         constructing_unit_Datapath_Middle_registers1_v_11_n66,
         constructing_unit_Datapath_Middle_registers1_v_11_n65,
         constructing_unit_Datapath_Middle_registers1_v_11_n64,
         constructing_unit_Datapath_Middle_registers1_v_11_n63,
         constructing_unit_Datapath_Middle_registers1_v_11_n62,
         constructing_unit_Datapath_Middle_registers1_v_11_n61,
         constructing_unit_Datapath_Middle_registers1_v_11_n60,
         constructing_unit_Datapath_Middle_registers1_v_11_n59,
         constructing_unit_Datapath_Middle_registers1_v_11_n58,
         constructing_unit_Datapath_Middle_registers1_v_11_n57,
         constructing_unit_Datapath_Middle_registers1_v_11_n56,
         constructing_unit_Datapath_Middle_registers1_v_11_n55,
         constructing_unit_Datapath_Middle_registers1_v_11_n54,
         constructing_unit_Datapath_Middle_registers1_v_11_n53,
         constructing_unit_Datapath_Middle_registers1_v_11_n52,
         constructing_unit_Datapath_Middle_registers1_v_11_n51,
         constructing_unit_Datapath_Middle_registers1_v_11_n50,
         constructing_unit_Datapath_Middle_registers1_v_11_n49,
         constructing_unit_Datapath_Middle_registers1_v_11_n48,
         constructing_unit_Datapath_Middle_registers1_v_11_n47,
         constructing_unit_Datapath_Middle_registers1_v_11_n46,
         constructing_unit_Datapath_Middle_registers1_v_11_n45,
         constructing_unit_Datapath_Middle_registers1_v_11_n44,
         constructing_unit_Datapath_Middle_registers1_v_11_n43,
         constructing_unit_Datapath_Middle_registers1_v_11_n42,
         constructing_unit_Datapath_Middle_registers1_v_11_n41,
         constructing_unit_Datapath_Middle_registers1_v_11_n40,
         constructing_unit_Datapath_Middle_registers1_v_11_n39,
         constructing_unit_Datapath_Middle_registers1_v_11_n38,
         constructing_unit_Datapath_Middle_registers1_v_11_n37,
         constructing_unit_Datapath_Middle_registers1_v_11_n36,
         constructing_unit_Datapath_Middle_registers1_v_11_n35,
         constructing_unit_Datapath_Middle_registers1_v_11_n33,
         constructing_unit_Datapath_Middle_registers1_v_12_n67,
         constructing_unit_Datapath_Middle_registers1_v_12_n66,
         constructing_unit_Datapath_Middle_registers1_v_12_n65,
         constructing_unit_Datapath_Middle_registers1_v_12_n64,
         constructing_unit_Datapath_Middle_registers1_v_12_n63,
         constructing_unit_Datapath_Middle_registers1_v_12_n62,
         constructing_unit_Datapath_Middle_registers1_v_12_n61,
         constructing_unit_Datapath_Middle_registers1_v_12_n60,
         constructing_unit_Datapath_Middle_registers1_v_12_n59,
         constructing_unit_Datapath_Middle_registers1_v_12_n58,
         constructing_unit_Datapath_Middle_registers1_v_12_n57,
         constructing_unit_Datapath_Middle_registers1_v_12_n56,
         constructing_unit_Datapath_Middle_registers1_v_12_n55,
         constructing_unit_Datapath_Middle_registers1_v_12_n54,
         constructing_unit_Datapath_Middle_registers1_v_12_n53,
         constructing_unit_Datapath_Middle_registers1_v_12_n52,
         constructing_unit_Datapath_Middle_registers1_v_12_n51,
         constructing_unit_Datapath_Middle_registers1_v_12_n50,
         constructing_unit_Datapath_Middle_registers1_v_12_n49,
         constructing_unit_Datapath_Middle_registers1_v_12_n48,
         constructing_unit_Datapath_Middle_registers1_v_12_n47,
         constructing_unit_Datapath_Middle_registers1_v_12_n46,
         constructing_unit_Datapath_Middle_registers1_v_12_n45,
         constructing_unit_Datapath_Middle_registers1_v_12_n44,
         constructing_unit_Datapath_Middle_registers1_v_12_n43,
         constructing_unit_Datapath_Middle_registers1_v_12_n42,
         constructing_unit_Datapath_Middle_registers1_v_12_n41,
         constructing_unit_Datapath_Middle_registers1_v_12_n40,
         constructing_unit_Datapath_Middle_registers1_v_12_n39,
         constructing_unit_Datapath_Middle_registers1_v_12_n38,
         constructing_unit_Datapath_Middle_registers1_v_12_n37,
         constructing_unit_Datapath_Middle_registers1_v_12_n36,
         constructing_unit_Datapath_Middle_registers1_v_12_n35,
         constructing_unit_Datapath_Middle_registers1_v_12_n33,
         constructing_unit_Datapath_Middle_registers1_v_13_n67,
         constructing_unit_Datapath_Middle_registers1_v_13_n66,
         constructing_unit_Datapath_Middle_registers1_v_13_n65,
         constructing_unit_Datapath_Middle_registers1_v_13_n64,
         constructing_unit_Datapath_Middle_registers1_v_13_n63,
         constructing_unit_Datapath_Middle_registers1_v_13_n62,
         constructing_unit_Datapath_Middle_registers1_v_13_n61,
         constructing_unit_Datapath_Middle_registers1_v_13_n60,
         constructing_unit_Datapath_Middle_registers1_v_13_n59,
         constructing_unit_Datapath_Middle_registers1_v_13_n58,
         constructing_unit_Datapath_Middle_registers1_v_13_n57,
         constructing_unit_Datapath_Middle_registers1_v_13_n56,
         constructing_unit_Datapath_Middle_registers1_v_13_n55,
         constructing_unit_Datapath_Middle_registers1_v_13_n54,
         constructing_unit_Datapath_Middle_registers1_v_13_n53,
         constructing_unit_Datapath_Middle_registers1_v_13_n52,
         constructing_unit_Datapath_Middle_registers1_v_13_n51,
         constructing_unit_Datapath_Middle_registers1_v_13_n50,
         constructing_unit_Datapath_Middle_registers1_v_13_n49,
         constructing_unit_Datapath_Middle_registers1_v_13_n48,
         constructing_unit_Datapath_Middle_registers1_v_13_n47,
         constructing_unit_Datapath_Middle_registers1_v_13_n46,
         constructing_unit_Datapath_Middle_registers1_v_13_n45,
         constructing_unit_Datapath_Middle_registers1_v_13_n44,
         constructing_unit_Datapath_Middle_registers1_v_13_n43,
         constructing_unit_Datapath_Middle_registers1_v_13_n42,
         constructing_unit_Datapath_Middle_registers1_v_13_n41,
         constructing_unit_Datapath_Middle_registers1_v_13_n40,
         constructing_unit_Datapath_Middle_registers1_v_13_n39,
         constructing_unit_Datapath_Middle_registers1_v_13_n38,
         constructing_unit_Datapath_Middle_registers1_v_13_n37,
         constructing_unit_Datapath_Middle_registers1_v_13_n36,
         constructing_unit_Datapath_Middle_registers1_v_13_n35,
         constructing_unit_Datapath_Middle_registers1_v_13_n33,
         constructing_unit_Datapath_Middle_registers2_v_3_n67,
         constructing_unit_Datapath_Middle_registers2_v_3_n66,
         constructing_unit_Datapath_Middle_registers2_v_3_n65,
         constructing_unit_Datapath_Middle_registers2_v_3_n64,
         constructing_unit_Datapath_Middle_registers2_v_3_n63,
         constructing_unit_Datapath_Middle_registers2_v_3_n62,
         constructing_unit_Datapath_Middle_registers2_v_3_n61,
         constructing_unit_Datapath_Middle_registers2_v_3_n60,
         constructing_unit_Datapath_Middle_registers2_v_3_n59,
         constructing_unit_Datapath_Middle_registers2_v_3_n58,
         constructing_unit_Datapath_Middle_registers2_v_3_n57,
         constructing_unit_Datapath_Middle_registers2_v_3_n56,
         constructing_unit_Datapath_Middle_registers2_v_3_n55,
         constructing_unit_Datapath_Middle_registers2_v_3_n54,
         constructing_unit_Datapath_Middle_registers2_v_3_n53,
         constructing_unit_Datapath_Middle_registers2_v_3_n52,
         constructing_unit_Datapath_Middle_registers2_v_3_n51,
         constructing_unit_Datapath_Middle_registers2_v_3_n50,
         constructing_unit_Datapath_Middle_registers2_v_3_n49,
         constructing_unit_Datapath_Middle_registers2_v_3_n48,
         constructing_unit_Datapath_Middle_registers2_v_3_n47,
         constructing_unit_Datapath_Middle_registers2_v_3_n46,
         constructing_unit_Datapath_Middle_registers2_v_3_n45,
         constructing_unit_Datapath_Middle_registers2_v_3_n44,
         constructing_unit_Datapath_Middle_registers2_v_3_n43,
         constructing_unit_Datapath_Middle_registers2_v_3_n42,
         constructing_unit_Datapath_Middle_registers2_v_3_n41,
         constructing_unit_Datapath_Middle_registers2_v_3_n40,
         constructing_unit_Datapath_Middle_registers2_v_3_n39,
         constructing_unit_Datapath_Middle_registers2_v_3_n38,
         constructing_unit_Datapath_Middle_registers2_v_3_n37,
         constructing_unit_Datapath_Middle_registers2_v_3_n36,
         constructing_unit_Datapath_Middle_registers2_v_3_n35,
         constructing_unit_Datapath_Middle_registers2_v_3_n33,
         constructing_unit_Datapath_Middle_registers2_v_4_n67,
         constructing_unit_Datapath_Middle_registers2_v_4_n66,
         constructing_unit_Datapath_Middle_registers2_v_4_n65,
         constructing_unit_Datapath_Middle_registers2_v_4_n64,
         constructing_unit_Datapath_Middle_registers2_v_4_n63,
         constructing_unit_Datapath_Middle_registers2_v_4_n62,
         constructing_unit_Datapath_Middle_registers2_v_4_n61,
         constructing_unit_Datapath_Middle_registers2_v_4_n60,
         constructing_unit_Datapath_Middle_registers2_v_4_n59,
         constructing_unit_Datapath_Middle_registers2_v_4_n58,
         constructing_unit_Datapath_Middle_registers2_v_4_n57,
         constructing_unit_Datapath_Middle_registers2_v_4_n56,
         constructing_unit_Datapath_Middle_registers2_v_4_n55,
         constructing_unit_Datapath_Middle_registers2_v_4_n54,
         constructing_unit_Datapath_Middle_registers2_v_4_n53,
         constructing_unit_Datapath_Middle_registers2_v_4_n52,
         constructing_unit_Datapath_Middle_registers2_v_4_n51,
         constructing_unit_Datapath_Middle_registers2_v_4_n50,
         constructing_unit_Datapath_Middle_registers2_v_4_n49,
         constructing_unit_Datapath_Middle_registers2_v_4_n48,
         constructing_unit_Datapath_Middle_registers2_v_4_n47,
         constructing_unit_Datapath_Middle_registers2_v_4_n46,
         constructing_unit_Datapath_Middle_registers2_v_4_n45,
         constructing_unit_Datapath_Middle_registers2_v_4_n44,
         constructing_unit_Datapath_Middle_registers2_v_4_n43,
         constructing_unit_Datapath_Middle_registers2_v_4_n42,
         constructing_unit_Datapath_Middle_registers2_v_4_n41,
         constructing_unit_Datapath_Middle_registers2_v_4_n40,
         constructing_unit_Datapath_Middle_registers2_v_4_n39,
         constructing_unit_Datapath_Middle_registers2_v_4_n38,
         constructing_unit_Datapath_Middle_registers2_v_4_n37,
         constructing_unit_Datapath_Middle_registers2_v_4_n36,
         constructing_unit_Datapath_Middle_registers2_v_4_n35,
         constructing_unit_Datapath_Middle_registers2_v_4_n33,
         constructing_unit_Datapath_Middle_registers2_v_5_n67,
         constructing_unit_Datapath_Middle_registers2_v_5_n66,
         constructing_unit_Datapath_Middle_registers2_v_5_n65,
         constructing_unit_Datapath_Middle_registers2_v_5_n64,
         constructing_unit_Datapath_Middle_registers2_v_5_n63,
         constructing_unit_Datapath_Middle_registers2_v_5_n62,
         constructing_unit_Datapath_Middle_registers2_v_5_n61,
         constructing_unit_Datapath_Middle_registers2_v_5_n60,
         constructing_unit_Datapath_Middle_registers2_v_5_n59,
         constructing_unit_Datapath_Middle_registers2_v_5_n58,
         constructing_unit_Datapath_Middle_registers2_v_5_n57,
         constructing_unit_Datapath_Middle_registers2_v_5_n56,
         constructing_unit_Datapath_Middle_registers2_v_5_n55,
         constructing_unit_Datapath_Middle_registers2_v_5_n54,
         constructing_unit_Datapath_Middle_registers2_v_5_n53,
         constructing_unit_Datapath_Middle_registers2_v_5_n52,
         constructing_unit_Datapath_Middle_registers2_v_5_n51,
         constructing_unit_Datapath_Middle_registers2_v_5_n50,
         constructing_unit_Datapath_Middle_registers2_v_5_n49,
         constructing_unit_Datapath_Middle_registers2_v_5_n48,
         constructing_unit_Datapath_Middle_registers2_v_5_n47,
         constructing_unit_Datapath_Middle_registers2_v_5_n46,
         constructing_unit_Datapath_Middle_registers2_v_5_n45,
         constructing_unit_Datapath_Middle_registers2_v_5_n44,
         constructing_unit_Datapath_Middle_registers2_v_5_n43,
         constructing_unit_Datapath_Middle_registers2_v_5_n42,
         constructing_unit_Datapath_Middle_registers2_v_5_n41,
         constructing_unit_Datapath_Middle_registers2_v_5_n40,
         constructing_unit_Datapath_Middle_registers2_v_5_n39,
         constructing_unit_Datapath_Middle_registers2_v_5_n38,
         constructing_unit_Datapath_Middle_registers2_v_5_n37,
         constructing_unit_Datapath_Middle_registers2_v_5_n36,
         constructing_unit_Datapath_Middle_registers2_v_5_n35,
         constructing_unit_Datapath_Middle_registers2_v_5_n33,
         constructing_unit_Datapath_Middle_registers2_v_6_n67,
         constructing_unit_Datapath_Middle_registers2_v_6_n66,
         constructing_unit_Datapath_Middle_registers2_v_6_n65,
         constructing_unit_Datapath_Middle_registers2_v_6_n64,
         constructing_unit_Datapath_Middle_registers2_v_6_n63,
         constructing_unit_Datapath_Middle_registers2_v_6_n62,
         constructing_unit_Datapath_Middle_registers2_v_6_n61,
         constructing_unit_Datapath_Middle_registers2_v_6_n60,
         constructing_unit_Datapath_Middle_registers2_v_6_n59,
         constructing_unit_Datapath_Middle_registers2_v_6_n58,
         constructing_unit_Datapath_Middle_registers2_v_6_n57,
         constructing_unit_Datapath_Middle_registers2_v_6_n56,
         constructing_unit_Datapath_Middle_registers2_v_6_n55,
         constructing_unit_Datapath_Middle_registers2_v_6_n54,
         constructing_unit_Datapath_Middle_registers2_v_6_n53,
         constructing_unit_Datapath_Middle_registers2_v_6_n52,
         constructing_unit_Datapath_Middle_registers2_v_6_n51,
         constructing_unit_Datapath_Middle_registers2_v_6_n50,
         constructing_unit_Datapath_Middle_registers2_v_6_n49,
         constructing_unit_Datapath_Middle_registers2_v_6_n48,
         constructing_unit_Datapath_Middle_registers2_v_6_n47,
         constructing_unit_Datapath_Middle_registers2_v_6_n46,
         constructing_unit_Datapath_Middle_registers2_v_6_n45,
         constructing_unit_Datapath_Middle_registers2_v_6_n44,
         constructing_unit_Datapath_Middle_registers2_v_6_n43,
         constructing_unit_Datapath_Middle_registers2_v_6_n42,
         constructing_unit_Datapath_Middle_registers2_v_6_n41,
         constructing_unit_Datapath_Middle_registers2_v_6_n40,
         constructing_unit_Datapath_Middle_registers2_v_6_n39,
         constructing_unit_Datapath_Middle_registers2_v_6_n38,
         constructing_unit_Datapath_Middle_registers2_v_6_n37,
         constructing_unit_Datapath_Middle_registers2_v_6_n36,
         constructing_unit_Datapath_Middle_registers2_v_6_n35,
         constructing_unit_Datapath_Middle_registers2_v_6_n33,
         constructing_unit_Datapath_Middle_registers2_v_7_n67,
         constructing_unit_Datapath_Middle_registers2_v_7_n66,
         constructing_unit_Datapath_Middle_registers2_v_7_n65,
         constructing_unit_Datapath_Middle_registers2_v_7_n64,
         constructing_unit_Datapath_Middle_registers2_v_7_n63,
         constructing_unit_Datapath_Middle_registers2_v_7_n62,
         constructing_unit_Datapath_Middle_registers2_v_7_n61,
         constructing_unit_Datapath_Middle_registers2_v_7_n60,
         constructing_unit_Datapath_Middle_registers2_v_7_n59,
         constructing_unit_Datapath_Middle_registers2_v_7_n58,
         constructing_unit_Datapath_Middle_registers2_v_7_n57,
         constructing_unit_Datapath_Middle_registers2_v_7_n56,
         constructing_unit_Datapath_Middle_registers2_v_7_n55,
         constructing_unit_Datapath_Middle_registers2_v_7_n54,
         constructing_unit_Datapath_Middle_registers2_v_7_n53,
         constructing_unit_Datapath_Middle_registers2_v_7_n52,
         constructing_unit_Datapath_Middle_registers2_v_7_n51,
         constructing_unit_Datapath_Middle_registers2_v_7_n50,
         constructing_unit_Datapath_Middle_registers2_v_7_n49,
         constructing_unit_Datapath_Middle_registers2_v_7_n48,
         constructing_unit_Datapath_Middle_registers2_v_7_n47,
         constructing_unit_Datapath_Middle_registers2_v_7_n46,
         constructing_unit_Datapath_Middle_registers2_v_7_n45,
         constructing_unit_Datapath_Middle_registers2_v_7_n44,
         constructing_unit_Datapath_Middle_registers2_v_7_n43,
         constructing_unit_Datapath_Middle_registers2_v_7_n42,
         constructing_unit_Datapath_Middle_registers2_v_7_n41,
         constructing_unit_Datapath_Middle_registers2_v_7_n40,
         constructing_unit_Datapath_Middle_registers2_v_7_n39,
         constructing_unit_Datapath_Middle_registers2_v_7_n38,
         constructing_unit_Datapath_Middle_registers2_v_7_n37,
         constructing_unit_Datapath_Middle_registers2_v_7_n36,
         constructing_unit_Datapath_Middle_registers2_v_7_n35,
         constructing_unit_Datapath_Middle_registers2_v_7_n33,
         constructing_unit_Datapath_Middle_registers2_v_8_n67,
         constructing_unit_Datapath_Middle_registers2_v_8_n66,
         constructing_unit_Datapath_Middle_registers2_v_8_n65,
         constructing_unit_Datapath_Middle_registers2_v_8_n64,
         constructing_unit_Datapath_Middle_registers2_v_8_n63,
         constructing_unit_Datapath_Middle_registers2_v_8_n62,
         constructing_unit_Datapath_Middle_registers2_v_8_n61,
         constructing_unit_Datapath_Middle_registers2_v_8_n60,
         constructing_unit_Datapath_Middle_registers2_v_8_n59,
         constructing_unit_Datapath_Middle_registers2_v_8_n58,
         constructing_unit_Datapath_Middle_registers2_v_8_n57,
         constructing_unit_Datapath_Middle_registers2_v_8_n56,
         constructing_unit_Datapath_Middle_registers2_v_8_n55,
         constructing_unit_Datapath_Middle_registers2_v_8_n54,
         constructing_unit_Datapath_Middle_registers2_v_8_n53,
         constructing_unit_Datapath_Middle_registers2_v_8_n52,
         constructing_unit_Datapath_Middle_registers2_v_8_n51,
         constructing_unit_Datapath_Middle_registers2_v_8_n50,
         constructing_unit_Datapath_Middle_registers2_v_8_n49,
         constructing_unit_Datapath_Middle_registers2_v_8_n48,
         constructing_unit_Datapath_Middle_registers2_v_8_n47,
         constructing_unit_Datapath_Middle_registers2_v_8_n46,
         constructing_unit_Datapath_Middle_registers2_v_8_n45,
         constructing_unit_Datapath_Middle_registers2_v_8_n44,
         constructing_unit_Datapath_Middle_registers2_v_8_n43,
         constructing_unit_Datapath_Middle_registers2_v_8_n42,
         constructing_unit_Datapath_Middle_registers2_v_8_n41,
         constructing_unit_Datapath_Middle_registers2_v_8_n40,
         constructing_unit_Datapath_Middle_registers2_v_8_n39,
         constructing_unit_Datapath_Middle_registers2_v_8_n38,
         constructing_unit_Datapath_Middle_registers2_v_8_n37,
         constructing_unit_Datapath_Middle_registers2_v_8_n36,
         constructing_unit_Datapath_Middle_registers2_v_8_n35,
         constructing_unit_Datapath_Middle_registers2_v_8_n33,
         constructing_unit_Datapath_Middle_registers2_v_9_n67,
         constructing_unit_Datapath_Middle_registers2_v_9_n66,
         constructing_unit_Datapath_Middle_registers2_v_9_n65,
         constructing_unit_Datapath_Middle_registers2_v_9_n64,
         constructing_unit_Datapath_Middle_registers2_v_9_n63,
         constructing_unit_Datapath_Middle_registers2_v_9_n62,
         constructing_unit_Datapath_Middle_registers2_v_9_n61,
         constructing_unit_Datapath_Middle_registers2_v_9_n60,
         constructing_unit_Datapath_Middle_registers2_v_9_n59,
         constructing_unit_Datapath_Middle_registers2_v_9_n58,
         constructing_unit_Datapath_Middle_registers2_v_9_n57,
         constructing_unit_Datapath_Middle_registers2_v_9_n56,
         constructing_unit_Datapath_Middle_registers2_v_9_n55,
         constructing_unit_Datapath_Middle_registers2_v_9_n54,
         constructing_unit_Datapath_Middle_registers2_v_9_n53,
         constructing_unit_Datapath_Middle_registers2_v_9_n52,
         constructing_unit_Datapath_Middle_registers2_v_9_n51,
         constructing_unit_Datapath_Middle_registers2_v_9_n50,
         constructing_unit_Datapath_Middle_registers2_v_9_n49,
         constructing_unit_Datapath_Middle_registers2_v_9_n48,
         constructing_unit_Datapath_Middle_registers2_v_9_n47,
         constructing_unit_Datapath_Middle_registers2_v_9_n46,
         constructing_unit_Datapath_Middle_registers2_v_9_n45,
         constructing_unit_Datapath_Middle_registers2_v_9_n44,
         constructing_unit_Datapath_Middle_registers2_v_9_n43,
         constructing_unit_Datapath_Middle_registers2_v_9_n42,
         constructing_unit_Datapath_Middle_registers2_v_9_n41,
         constructing_unit_Datapath_Middle_registers2_v_9_n40,
         constructing_unit_Datapath_Middle_registers2_v_9_n39,
         constructing_unit_Datapath_Middle_registers2_v_9_n38,
         constructing_unit_Datapath_Middle_registers2_v_9_n37,
         constructing_unit_Datapath_Middle_registers2_v_9_n36,
         constructing_unit_Datapath_Middle_registers2_v_9_n35,
         constructing_unit_Datapath_Middle_registers2_v_9_n33,
         constructing_unit_Datapath_Middle_registers2_v_10_n67,
         constructing_unit_Datapath_Middle_registers2_v_10_n66,
         constructing_unit_Datapath_Middle_registers2_v_10_n65,
         constructing_unit_Datapath_Middle_registers2_v_10_n64,
         constructing_unit_Datapath_Middle_registers2_v_10_n63,
         constructing_unit_Datapath_Middle_registers2_v_10_n62,
         constructing_unit_Datapath_Middle_registers2_v_10_n61,
         constructing_unit_Datapath_Middle_registers2_v_10_n60,
         constructing_unit_Datapath_Middle_registers2_v_10_n59,
         constructing_unit_Datapath_Middle_registers2_v_10_n58,
         constructing_unit_Datapath_Middle_registers2_v_10_n57,
         constructing_unit_Datapath_Middle_registers2_v_10_n56,
         constructing_unit_Datapath_Middle_registers2_v_10_n55,
         constructing_unit_Datapath_Middle_registers2_v_10_n54,
         constructing_unit_Datapath_Middle_registers2_v_10_n53,
         constructing_unit_Datapath_Middle_registers2_v_10_n52,
         constructing_unit_Datapath_Middle_registers2_v_10_n51,
         constructing_unit_Datapath_Middle_registers2_v_10_n50,
         constructing_unit_Datapath_Middle_registers2_v_10_n49,
         constructing_unit_Datapath_Middle_registers2_v_10_n48,
         constructing_unit_Datapath_Middle_registers2_v_10_n47,
         constructing_unit_Datapath_Middle_registers2_v_10_n46,
         constructing_unit_Datapath_Middle_registers2_v_10_n45,
         constructing_unit_Datapath_Middle_registers2_v_10_n44,
         constructing_unit_Datapath_Middle_registers2_v_10_n43,
         constructing_unit_Datapath_Middle_registers2_v_10_n42,
         constructing_unit_Datapath_Middle_registers2_v_10_n41,
         constructing_unit_Datapath_Middle_registers2_v_10_n40,
         constructing_unit_Datapath_Middle_registers2_v_10_n39,
         constructing_unit_Datapath_Middle_registers2_v_10_n38,
         constructing_unit_Datapath_Middle_registers2_v_10_n37,
         constructing_unit_Datapath_Middle_registers2_v_10_n36,
         constructing_unit_Datapath_Middle_registers2_v_10_n35,
         constructing_unit_Datapath_Middle_registers2_v_10_n33,
         constructing_unit_Datapath_Middle_registers2_v_11_n67,
         constructing_unit_Datapath_Middle_registers2_v_11_n66,
         constructing_unit_Datapath_Middle_registers2_v_11_n65,
         constructing_unit_Datapath_Middle_registers2_v_11_n64,
         constructing_unit_Datapath_Middle_registers2_v_11_n63,
         constructing_unit_Datapath_Middle_registers2_v_11_n62,
         constructing_unit_Datapath_Middle_registers2_v_11_n61,
         constructing_unit_Datapath_Middle_registers2_v_11_n60,
         constructing_unit_Datapath_Middle_registers2_v_11_n59,
         constructing_unit_Datapath_Middle_registers2_v_11_n58,
         constructing_unit_Datapath_Middle_registers2_v_11_n57,
         constructing_unit_Datapath_Middle_registers2_v_11_n56,
         constructing_unit_Datapath_Middle_registers2_v_11_n55,
         constructing_unit_Datapath_Middle_registers2_v_11_n54,
         constructing_unit_Datapath_Middle_registers2_v_11_n53,
         constructing_unit_Datapath_Middle_registers2_v_11_n52,
         constructing_unit_Datapath_Middle_registers2_v_11_n51,
         constructing_unit_Datapath_Middle_registers2_v_11_n50,
         constructing_unit_Datapath_Middle_registers2_v_11_n49,
         constructing_unit_Datapath_Middle_registers2_v_11_n48,
         constructing_unit_Datapath_Middle_registers2_v_11_n47,
         constructing_unit_Datapath_Middle_registers2_v_11_n46,
         constructing_unit_Datapath_Middle_registers2_v_11_n45,
         constructing_unit_Datapath_Middle_registers2_v_11_n44,
         constructing_unit_Datapath_Middle_registers2_v_11_n43,
         constructing_unit_Datapath_Middle_registers2_v_11_n42,
         constructing_unit_Datapath_Middle_registers2_v_11_n41,
         constructing_unit_Datapath_Middle_registers2_v_11_n40,
         constructing_unit_Datapath_Middle_registers2_v_11_n39,
         constructing_unit_Datapath_Middle_registers2_v_11_n38,
         constructing_unit_Datapath_Middle_registers2_v_11_n37,
         constructing_unit_Datapath_Middle_registers2_v_11_n36,
         constructing_unit_Datapath_Middle_registers2_v_11_n35,
         constructing_unit_Datapath_Middle_registers2_v_11_n33,
         constructing_unit_Datapath_Middle_registers2_v_12_n67,
         constructing_unit_Datapath_Middle_registers2_v_12_n66,
         constructing_unit_Datapath_Middle_registers2_v_12_n65,
         constructing_unit_Datapath_Middle_registers2_v_12_n64,
         constructing_unit_Datapath_Middle_registers2_v_12_n63,
         constructing_unit_Datapath_Middle_registers2_v_12_n62,
         constructing_unit_Datapath_Middle_registers2_v_12_n61,
         constructing_unit_Datapath_Middle_registers2_v_12_n60,
         constructing_unit_Datapath_Middle_registers2_v_12_n59,
         constructing_unit_Datapath_Middle_registers2_v_12_n58,
         constructing_unit_Datapath_Middle_registers2_v_12_n57,
         constructing_unit_Datapath_Middle_registers2_v_12_n56,
         constructing_unit_Datapath_Middle_registers2_v_12_n55,
         constructing_unit_Datapath_Middle_registers2_v_12_n54,
         constructing_unit_Datapath_Middle_registers2_v_12_n53,
         constructing_unit_Datapath_Middle_registers2_v_12_n52,
         constructing_unit_Datapath_Middle_registers2_v_12_n51,
         constructing_unit_Datapath_Middle_registers2_v_12_n50,
         constructing_unit_Datapath_Middle_registers2_v_12_n49,
         constructing_unit_Datapath_Middle_registers2_v_12_n48,
         constructing_unit_Datapath_Middle_registers2_v_12_n47,
         constructing_unit_Datapath_Middle_registers2_v_12_n46,
         constructing_unit_Datapath_Middle_registers2_v_12_n45,
         constructing_unit_Datapath_Middle_registers2_v_12_n44,
         constructing_unit_Datapath_Middle_registers2_v_12_n43,
         constructing_unit_Datapath_Middle_registers2_v_12_n42,
         constructing_unit_Datapath_Middle_registers2_v_12_n41,
         constructing_unit_Datapath_Middle_registers2_v_12_n40,
         constructing_unit_Datapath_Middle_registers2_v_12_n39,
         constructing_unit_Datapath_Middle_registers2_v_12_n38,
         constructing_unit_Datapath_Middle_registers2_v_12_n37,
         constructing_unit_Datapath_Middle_registers2_v_12_n36,
         constructing_unit_Datapath_Middle_registers2_v_12_n35,
         constructing_unit_Datapath_Middle_registers2_v_12_n33,
         constructing_unit_Datapath_Middle_registers2_v_13_n67,
         constructing_unit_Datapath_Middle_registers2_v_13_n66,
         constructing_unit_Datapath_Middle_registers2_v_13_n65,
         constructing_unit_Datapath_Middle_registers2_v_13_n64,
         constructing_unit_Datapath_Middle_registers2_v_13_n63,
         constructing_unit_Datapath_Middle_registers2_v_13_n62,
         constructing_unit_Datapath_Middle_registers2_v_13_n61,
         constructing_unit_Datapath_Middle_registers2_v_13_n60,
         constructing_unit_Datapath_Middle_registers2_v_13_n59,
         constructing_unit_Datapath_Middle_registers2_v_13_n58,
         constructing_unit_Datapath_Middle_registers2_v_13_n57,
         constructing_unit_Datapath_Middle_registers2_v_13_n56,
         constructing_unit_Datapath_Middle_registers2_v_13_n55,
         constructing_unit_Datapath_Middle_registers2_v_13_n54,
         constructing_unit_Datapath_Middle_registers2_v_13_n53,
         constructing_unit_Datapath_Middle_registers2_v_13_n52,
         constructing_unit_Datapath_Middle_registers2_v_13_n51,
         constructing_unit_Datapath_Middle_registers2_v_13_n50,
         constructing_unit_Datapath_Middle_registers2_v_13_n49,
         constructing_unit_Datapath_Middle_registers2_v_13_n48,
         constructing_unit_Datapath_Middle_registers2_v_13_n47,
         constructing_unit_Datapath_Middle_registers2_v_13_n46,
         constructing_unit_Datapath_Middle_registers2_v_13_n45,
         constructing_unit_Datapath_Middle_registers2_v_13_n44,
         constructing_unit_Datapath_Middle_registers2_v_13_n43,
         constructing_unit_Datapath_Middle_registers2_v_13_n42,
         constructing_unit_Datapath_Middle_registers2_v_13_n41,
         constructing_unit_Datapath_Middle_registers2_v_13_n40,
         constructing_unit_Datapath_Middle_registers2_v_13_n39,
         constructing_unit_Datapath_Middle_registers2_v_13_n38,
         constructing_unit_Datapath_Middle_registers2_v_13_n37,
         constructing_unit_Datapath_Middle_registers2_v_13_n36,
         constructing_unit_Datapath_Middle_registers2_v_13_n35,
         constructing_unit_Datapath_Middle_registers2_v_13_n33,
         constructing_unit_Datapath_Last_register0_v_n69,
         constructing_unit_Datapath_Last_register0_v_n68,
         constructing_unit_Datapath_Last_register0_v_n67,
         constructing_unit_Datapath_Last_register0_v_n66,
         constructing_unit_Datapath_Last_register0_v_n65,
         constructing_unit_Datapath_Last_register0_v_n64,
         constructing_unit_Datapath_Last_register0_v_n63,
         constructing_unit_Datapath_Last_register0_v_n62,
         constructing_unit_Datapath_Last_register0_v_n61,
         constructing_unit_Datapath_Last_register0_v_n60,
         constructing_unit_Datapath_Last_register0_v_n59,
         constructing_unit_Datapath_Last_register0_v_n58,
         constructing_unit_Datapath_Last_register0_v_n57,
         constructing_unit_Datapath_Last_register0_v_n56,
         constructing_unit_Datapath_Last_register0_v_n55,
         constructing_unit_Datapath_Last_register0_v_n54,
         constructing_unit_Datapath_Last_register0_v_n53,
         constructing_unit_Datapath_Last_register0_v_n52,
         constructing_unit_Datapath_Last_register0_v_n51,
         constructing_unit_Datapath_Last_register0_v_n50,
         constructing_unit_Datapath_Last_register0_v_n49,
         constructing_unit_Datapath_Last_register0_v_n48,
         constructing_unit_Datapath_Last_register0_v_n47,
         constructing_unit_Datapath_Last_register0_v_n46,
         constructing_unit_Datapath_Last_register0_v_n45,
         constructing_unit_Datapath_Last_register0_v_n44,
         constructing_unit_Datapath_Last_register0_v_n43,
         constructing_unit_Datapath_Last_register0_v_n42,
         constructing_unit_Datapath_Last_register0_v_n41,
         constructing_unit_Datapath_Last_register0_v_n40,
         constructing_unit_Datapath_Last_register0_v_n39,
         constructing_unit_Datapath_Last_register0_v_n38,
         constructing_unit_Datapath_Last_register0_v_n37,
         constructing_unit_Datapath_Last_register0_v_n36,
         constructing_unit_Datapath_Last_register0_v_n35,
         constructing_unit_Datapath_Last_register0_v_n33,
         constructing_unit_Datapath_Last_register1_v_n69,
         constructing_unit_Datapath_Last_register1_v_n68,
         constructing_unit_Datapath_Last_register1_v_n67,
         constructing_unit_Datapath_Last_register1_v_n66,
         constructing_unit_Datapath_Last_register1_v_n65,
         constructing_unit_Datapath_Last_register1_v_n64,
         constructing_unit_Datapath_Last_register1_v_n63,
         constructing_unit_Datapath_Last_register1_v_n62,
         constructing_unit_Datapath_Last_register1_v_n61,
         constructing_unit_Datapath_Last_register1_v_n60,
         constructing_unit_Datapath_Last_register1_v_n59,
         constructing_unit_Datapath_Last_register1_v_n58,
         constructing_unit_Datapath_Last_register1_v_n57,
         constructing_unit_Datapath_Last_register1_v_n56,
         constructing_unit_Datapath_Last_register1_v_n55,
         constructing_unit_Datapath_Last_register1_v_n54,
         constructing_unit_Datapath_Last_register1_v_n53,
         constructing_unit_Datapath_Last_register1_v_n52,
         constructing_unit_Datapath_Last_register1_v_n51,
         constructing_unit_Datapath_Last_register1_v_n50,
         constructing_unit_Datapath_Last_register1_v_n49,
         constructing_unit_Datapath_Last_register1_v_n48,
         constructing_unit_Datapath_Last_register1_v_n47,
         constructing_unit_Datapath_Last_register1_v_n46,
         constructing_unit_Datapath_Last_register1_v_n45,
         constructing_unit_Datapath_Last_register1_v_n44,
         constructing_unit_Datapath_Last_register1_v_n43,
         constructing_unit_Datapath_Last_register1_v_n42,
         constructing_unit_Datapath_Last_register1_v_n41,
         constructing_unit_Datapath_Last_register1_v_n40,
         constructing_unit_Datapath_Last_register1_v_n39,
         constructing_unit_Datapath_Last_register1_v_n38,
         constructing_unit_Datapath_Last_register1_v_n37,
         constructing_unit_Datapath_Last_register1_v_n36,
         constructing_unit_Datapath_Last_register1_v_n35,
         constructing_unit_Datapath_Last_register1_v_n33,
         constructing_unit_Datapath_Last_register2_v_n69,
         constructing_unit_Datapath_Last_register2_v_n68,
         constructing_unit_Datapath_Last_register2_v_n67,
         constructing_unit_Datapath_Last_register2_v_n66,
         constructing_unit_Datapath_Last_register2_v_n65,
         constructing_unit_Datapath_Last_register2_v_n64,
         constructing_unit_Datapath_Last_register2_v_n63,
         constructing_unit_Datapath_Last_register2_v_n62,
         constructing_unit_Datapath_Last_register2_v_n61,
         constructing_unit_Datapath_Last_register2_v_n60,
         constructing_unit_Datapath_Last_register2_v_n59,
         constructing_unit_Datapath_Last_register2_v_n58,
         constructing_unit_Datapath_Last_register2_v_n57,
         constructing_unit_Datapath_Last_register2_v_n56,
         constructing_unit_Datapath_Last_register2_v_n55,
         constructing_unit_Datapath_Last_register2_v_n54,
         constructing_unit_Datapath_Last_register2_v_n53,
         constructing_unit_Datapath_Last_register2_v_n52,
         constructing_unit_Datapath_Last_register2_v_n51,
         constructing_unit_Datapath_Last_register2_v_n50,
         constructing_unit_Datapath_Last_register2_v_n49,
         constructing_unit_Datapath_Last_register2_v_n48,
         constructing_unit_Datapath_Last_register2_v_n47,
         constructing_unit_Datapath_Last_register2_v_n46,
         constructing_unit_Datapath_Last_register2_v_n45,
         constructing_unit_Datapath_Last_register2_v_n44,
         constructing_unit_Datapath_Last_register2_v_n43,
         constructing_unit_Datapath_Last_register2_v_n42,
         constructing_unit_Datapath_Last_register2_v_n41,
         constructing_unit_Datapath_Last_register2_v_n40,
         constructing_unit_Datapath_Last_register2_v_n39,
         constructing_unit_Datapath_Last_register2_v_n38,
         constructing_unit_Datapath_Last_register2_v_n37,
         constructing_unit_Datapath_Last_register2_v_n36,
         constructing_unit_Datapath_Last_register2_v_n35,
         constructing_unit_Datapath_Last_register2_v_n33,
         constructing_unit_Datapath_FaS_registers0_h_1_n67,
         constructing_unit_Datapath_FaS_registers0_h_1_n66,
         constructing_unit_Datapath_FaS_registers0_h_1_n65,
         constructing_unit_Datapath_FaS_registers0_h_1_n64,
         constructing_unit_Datapath_FaS_registers0_h_1_n63,
         constructing_unit_Datapath_FaS_registers0_h_1_n62,
         constructing_unit_Datapath_FaS_registers0_h_1_n61,
         constructing_unit_Datapath_FaS_registers0_h_1_n60,
         constructing_unit_Datapath_FaS_registers0_h_1_n59,
         constructing_unit_Datapath_FaS_registers0_h_1_n58,
         constructing_unit_Datapath_FaS_registers0_h_1_n57,
         constructing_unit_Datapath_FaS_registers0_h_1_n56,
         constructing_unit_Datapath_FaS_registers0_h_1_n55,
         constructing_unit_Datapath_FaS_registers0_h_1_n54,
         constructing_unit_Datapath_FaS_registers0_h_1_n53,
         constructing_unit_Datapath_FaS_registers0_h_1_n52,
         constructing_unit_Datapath_FaS_registers0_h_1_n51,
         constructing_unit_Datapath_FaS_registers0_h_1_n50,
         constructing_unit_Datapath_FaS_registers0_h_1_n49,
         constructing_unit_Datapath_FaS_registers0_h_1_n48,
         constructing_unit_Datapath_FaS_registers0_h_1_n47,
         constructing_unit_Datapath_FaS_registers0_h_1_n46,
         constructing_unit_Datapath_FaS_registers0_h_1_n45,
         constructing_unit_Datapath_FaS_registers0_h_1_n44,
         constructing_unit_Datapath_FaS_registers0_h_1_n43,
         constructing_unit_Datapath_FaS_registers0_h_1_n42,
         constructing_unit_Datapath_FaS_registers0_h_1_n41,
         constructing_unit_Datapath_FaS_registers0_h_1_n40,
         constructing_unit_Datapath_FaS_registers0_h_1_n39,
         constructing_unit_Datapath_FaS_registers0_h_1_n38,
         constructing_unit_Datapath_FaS_registers0_h_1_n37,
         constructing_unit_Datapath_FaS_registers0_h_1_n36,
         constructing_unit_Datapath_FaS_registers0_h_1_n35,
         constructing_unit_Datapath_FaS_registers0_h_1_n33,
         constructing_unit_Datapath_FaS_registers0_h_2_n67,
         constructing_unit_Datapath_FaS_registers0_h_2_n66,
         constructing_unit_Datapath_FaS_registers0_h_2_n65,
         constructing_unit_Datapath_FaS_registers0_h_2_n64,
         constructing_unit_Datapath_FaS_registers0_h_2_n63,
         constructing_unit_Datapath_FaS_registers0_h_2_n62,
         constructing_unit_Datapath_FaS_registers0_h_2_n61,
         constructing_unit_Datapath_FaS_registers0_h_2_n60,
         constructing_unit_Datapath_FaS_registers0_h_2_n59,
         constructing_unit_Datapath_FaS_registers0_h_2_n58,
         constructing_unit_Datapath_FaS_registers0_h_2_n57,
         constructing_unit_Datapath_FaS_registers0_h_2_n56,
         constructing_unit_Datapath_FaS_registers0_h_2_n55,
         constructing_unit_Datapath_FaS_registers0_h_2_n54,
         constructing_unit_Datapath_FaS_registers0_h_2_n53,
         constructing_unit_Datapath_FaS_registers0_h_2_n52,
         constructing_unit_Datapath_FaS_registers0_h_2_n51,
         constructing_unit_Datapath_FaS_registers0_h_2_n50,
         constructing_unit_Datapath_FaS_registers0_h_2_n49,
         constructing_unit_Datapath_FaS_registers0_h_2_n48,
         constructing_unit_Datapath_FaS_registers0_h_2_n47,
         constructing_unit_Datapath_FaS_registers0_h_2_n46,
         constructing_unit_Datapath_FaS_registers0_h_2_n45,
         constructing_unit_Datapath_FaS_registers0_h_2_n44,
         constructing_unit_Datapath_FaS_registers0_h_2_n43,
         constructing_unit_Datapath_FaS_registers0_h_2_n42,
         constructing_unit_Datapath_FaS_registers0_h_2_n41,
         constructing_unit_Datapath_FaS_registers0_h_2_n40,
         constructing_unit_Datapath_FaS_registers0_h_2_n39,
         constructing_unit_Datapath_FaS_registers0_h_2_n38,
         constructing_unit_Datapath_FaS_registers0_h_2_n37,
         constructing_unit_Datapath_FaS_registers0_h_2_n36,
         constructing_unit_Datapath_FaS_registers0_h_2_n35,
         constructing_unit_Datapath_FaS_registers0_h_2_n33,
         constructing_unit_Datapath_FaS_registers1_h_1_n67,
         constructing_unit_Datapath_FaS_registers1_h_1_n66,
         constructing_unit_Datapath_FaS_registers1_h_1_n65,
         constructing_unit_Datapath_FaS_registers1_h_1_n64,
         constructing_unit_Datapath_FaS_registers1_h_1_n63,
         constructing_unit_Datapath_FaS_registers1_h_1_n62,
         constructing_unit_Datapath_FaS_registers1_h_1_n61,
         constructing_unit_Datapath_FaS_registers1_h_1_n60,
         constructing_unit_Datapath_FaS_registers1_h_1_n59,
         constructing_unit_Datapath_FaS_registers1_h_1_n58,
         constructing_unit_Datapath_FaS_registers1_h_1_n57,
         constructing_unit_Datapath_FaS_registers1_h_1_n56,
         constructing_unit_Datapath_FaS_registers1_h_1_n55,
         constructing_unit_Datapath_FaS_registers1_h_1_n54,
         constructing_unit_Datapath_FaS_registers1_h_1_n53,
         constructing_unit_Datapath_FaS_registers1_h_1_n52,
         constructing_unit_Datapath_FaS_registers1_h_1_n51,
         constructing_unit_Datapath_FaS_registers1_h_1_n50,
         constructing_unit_Datapath_FaS_registers1_h_1_n49,
         constructing_unit_Datapath_FaS_registers1_h_1_n48,
         constructing_unit_Datapath_FaS_registers1_h_1_n47,
         constructing_unit_Datapath_FaS_registers1_h_1_n46,
         constructing_unit_Datapath_FaS_registers1_h_1_n45,
         constructing_unit_Datapath_FaS_registers1_h_1_n44,
         constructing_unit_Datapath_FaS_registers1_h_1_n43,
         constructing_unit_Datapath_FaS_registers1_h_1_n42,
         constructing_unit_Datapath_FaS_registers1_h_1_n41,
         constructing_unit_Datapath_FaS_registers1_h_1_n40,
         constructing_unit_Datapath_FaS_registers1_h_1_n39,
         constructing_unit_Datapath_FaS_registers1_h_1_n38,
         constructing_unit_Datapath_FaS_registers1_h_1_n37,
         constructing_unit_Datapath_FaS_registers1_h_1_n36,
         constructing_unit_Datapath_FaS_registers1_h_1_n35,
         constructing_unit_Datapath_FaS_registers1_h_1_n33,
         constructing_unit_Datapath_FaS_registers1_h_2_n67,
         constructing_unit_Datapath_FaS_registers1_h_2_n66,
         constructing_unit_Datapath_FaS_registers1_h_2_n65,
         constructing_unit_Datapath_FaS_registers1_h_2_n64,
         constructing_unit_Datapath_FaS_registers1_h_2_n63,
         constructing_unit_Datapath_FaS_registers1_h_2_n62,
         constructing_unit_Datapath_FaS_registers1_h_2_n61,
         constructing_unit_Datapath_FaS_registers1_h_2_n60,
         constructing_unit_Datapath_FaS_registers1_h_2_n59,
         constructing_unit_Datapath_FaS_registers1_h_2_n58,
         constructing_unit_Datapath_FaS_registers1_h_2_n57,
         constructing_unit_Datapath_FaS_registers1_h_2_n56,
         constructing_unit_Datapath_FaS_registers1_h_2_n55,
         constructing_unit_Datapath_FaS_registers1_h_2_n54,
         constructing_unit_Datapath_FaS_registers1_h_2_n53,
         constructing_unit_Datapath_FaS_registers1_h_2_n52,
         constructing_unit_Datapath_FaS_registers1_h_2_n51,
         constructing_unit_Datapath_FaS_registers1_h_2_n50,
         constructing_unit_Datapath_FaS_registers1_h_2_n49,
         constructing_unit_Datapath_FaS_registers1_h_2_n48,
         constructing_unit_Datapath_FaS_registers1_h_2_n47,
         constructing_unit_Datapath_FaS_registers1_h_2_n46,
         constructing_unit_Datapath_FaS_registers1_h_2_n45,
         constructing_unit_Datapath_FaS_registers1_h_2_n44,
         constructing_unit_Datapath_FaS_registers1_h_2_n43,
         constructing_unit_Datapath_FaS_registers1_h_2_n42,
         constructing_unit_Datapath_FaS_registers1_h_2_n41,
         constructing_unit_Datapath_FaS_registers1_h_2_n40,
         constructing_unit_Datapath_FaS_registers1_h_2_n39,
         constructing_unit_Datapath_FaS_registers1_h_2_n38,
         constructing_unit_Datapath_FaS_registers1_h_2_n37,
         constructing_unit_Datapath_FaS_registers1_h_2_n36,
         constructing_unit_Datapath_FaS_registers1_h_2_n35,
         constructing_unit_Datapath_FaS_registers1_h_2_n33,
         constructing_unit_Datapath_FaS_registers2_h_1_n67,
         constructing_unit_Datapath_FaS_registers2_h_1_n66,
         constructing_unit_Datapath_FaS_registers2_h_1_n65,
         constructing_unit_Datapath_FaS_registers2_h_1_n64,
         constructing_unit_Datapath_FaS_registers2_h_1_n63,
         constructing_unit_Datapath_FaS_registers2_h_1_n62,
         constructing_unit_Datapath_FaS_registers2_h_1_n61,
         constructing_unit_Datapath_FaS_registers2_h_1_n60,
         constructing_unit_Datapath_FaS_registers2_h_1_n59,
         constructing_unit_Datapath_FaS_registers2_h_1_n58,
         constructing_unit_Datapath_FaS_registers2_h_1_n57,
         constructing_unit_Datapath_FaS_registers2_h_1_n56,
         constructing_unit_Datapath_FaS_registers2_h_1_n55,
         constructing_unit_Datapath_FaS_registers2_h_1_n54,
         constructing_unit_Datapath_FaS_registers2_h_1_n53,
         constructing_unit_Datapath_FaS_registers2_h_1_n52,
         constructing_unit_Datapath_FaS_registers2_h_1_n51,
         constructing_unit_Datapath_FaS_registers2_h_1_n50,
         constructing_unit_Datapath_FaS_registers2_h_1_n49,
         constructing_unit_Datapath_FaS_registers2_h_1_n48,
         constructing_unit_Datapath_FaS_registers2_h_1_n47,
         constructing_unit_Datapath_FaS_registers2_h_1_n46,
         constructing_unit_Datapath_FaS_registers2_h_1_n45,
         constructing_unit_Datapath_FaS_registers2_h_1_n44,
         constructing_unit_Datapath_FaS_registers2_h_1_n43,
         constructing_unit_Datapath_FaS_registers2_h_1_n42,
         constructing_unit_Datapath_FaS_registers2_h_1_n41,
         constructing_unit_Datapath_FaS_registers2_h_1_n40,
         constructing_unit_Datapath_FaS_registers2_h_1_n39,
         constructing_unit_Datapath_FaS_registers2_h_1_n38,
         constructing_unit_Datapath_FaS_registers2_h_1_n37,
         constructing_unit_Datapath_FaS_registers2_h_1_n36,
         constructing_unit_Datapath_FaS_registers2_h_1_n35,
         constructing_unit_Datapath_FaS_registers2_h_1_n33,
         constructing_unit_Datapath_FaS_registers2_h_2_n67,
         constructing_unit_Datapath_FaS_registers2_h_2_n66,
         constructing_unit_Datapath_FaS_registers2_h_2_n65,
         constructing_unit_Datapath_FaS_registers2_h_2_n64,
         constructing_unit_Datapath_FaS_registers2_h_2_n63,
         constructing_unit_Datapath_FaS_registers2_h_2_n62,
         constructing_unit_Datapath_FaS_registers2_h_2_n61,
         constructing_unit_Datapath_FaS_registers2_h_2_n60,
         constructing_unit_Datapath_FaS_registers2_h_2_n59,
         constructing_unit_Datapath_FaS_registers2_h_2_n58,
         constructing_unit_Datapath_FaS_registers2_h_2_n57,
         constructing_unit_Datapath_FaS_registers2_h_2_n56,
         constructing_unit_Datapath_FaS_registers2_h_2_n55,
         constructing_unit_Datapath_FaS_registers2_h_2_n54,
         constructing_unit_Datapath_FaS_registers2_h_2_n53,
         constructing_unit_Datapath_FaS_registers2_h_2_n52,
         constructing_unit_Datapath_FaS_registers2_h_2_n51,
         constructing_unit_Datapath_FaS_registers2_h_2_n50,
         constructing_unit_Datapath_FaS_registers2_h_2_n49,
         constructing_unit_Datapath_FaS_registers2_h_2_n48,
         constructing_unit_Datapath_FaS_registers2_h_2_n47,
         constructing_unit_Datapath_FaS_registers2_h_2_n46,
         constructing_unit_Datapath_FaS_registers2_h_2_n45,
         constructing_unit_Datapath_FaS_registers2_h_2_n44,
         constructing_unit_Datapath_FaS_registers2_h_2_n43,
         constructing_unit_Datapath_FaS_registers2_h_2_n42,
         constructing_unit_Datapath_FaS_registers2_h_2_n41,
         constructing_unit_Datapath_FaS_registers2_h_2_n40,
         constructing_unit_Datapath_FaS_registers2_h_2_n39,
         constructing_unit_Datapath_FaS_registers2_h_2_n38,
         constructing_unit_Datapath_FaS_registers2_h_2_n37,
         constructing_unit_Datapath_FaS_registers2_h_2_n36,
         constructing_unit_Datapath_FaS_registers2_h_2_n35,
         constructing_unit_Datapath_FaS_registers2_h_2_n33,
         constructing_unit_Datapath_Middle_registers0_h_3_n67,
         constructing_unit_Datapath_Middle_registers0_h_3_n66,
         constructing_unit_Datapath_Middle_registers0_h_3_n65,
         constructing_unit_Datapath_Middle_registers0_h_3_n64,
         constructing_unit_Datapath_Middle_registers0_h_3_n63,
         constructing_unit_Datapath_Middle_registers0_h_3_n62,
         constructing_unit_Datapath_Middle_registers0_h_3_n61,
         constructing_unit_Datapath_Middle_registers0_h_3_n60,
         constructing_unit_Datapath_Middle_registers0_h_3_n59,
         constructing_unit_Datapath_Middle_registers0_h_3_n58,
         constructing_unit_Datapath_Middle_registers0_h_3_n57,
         constructing_unit_Datapath_Middle_registers0_h_3_n56,
         constructing_unit_Datapath_Middle_registers0_h_3_n55,
         constructing_unit_Datapath_Middle_registers0_h_3_n54,
         constructing_unit_Datapath_Middle_registers0_h_3_n53,
         constructing_unit_Datapath_Middle_registers0_h_3_n52,
         constructing_unit_Datapath_Middle_registers0_h_3_n51,
         constructing_unit_Datapath_Middle_registers0_h_3_n50,
         constructing_unit_Datapath_Middle_registers0_h_3_n49,
         constructing_unit_Datapath_Middle_registers0_h_3_n48,
         constructing_unit_Datapath_Middle_registers0_h_3_n47,
         constructing_unit_Datapath_Middle_registers0_h_3_n46,
         constructing_unit_Datapath_Middle_registers0_h_3_n45,
         constructing_unit_Datapath_Middle_registers0_h_3_n44,
         constructing_unit_Datapath_Middle_registers0_h_3_n43,
         constructing_unit_Datapath_Middle_registers0_h_3_n42,
         constructing_unit_Datapath_Middle_registers0_h_3_n41,
         constructing_unit_Datapath_Middle_registers0_h_3_n40,
         constructing_unit_Datapath_Middle_registers0_h_3_n39,
         constructing_unit_Datapath_Middle_registers0_h_3_n38,
         constructing_unit_Datapath_Middle_registers0_h_3_n37,
         constructing_unit_Datapath_Middle_registers0_h_3_n36,
         constructing_unit_Datapath_Middle_registers0_h_3_n35,
         constructing_unit_Datapath_Middle_registers0_h_3_n33,
         constructing_unit_Datapath_Middle_registers0_h_4_n67,
         constructing_unit_Datapath_Middle_registers0_h_4_n66,
         constructing_unit_Datapath_Middle_registers0_h_4_n65,
         constructing_unit_Datapath_Middle_registers0_h_4_n64,
         constructing_unit_Datapath_Middle_registers0_h_4_n63,
         constructing_unit_Datapath_Middle_registers0_h_4_n62,
         constructing_unit_Datapath_Middle_registers0_h_4_n61,
         constructing_unit_Datapath_Middle_registers0_h_4_n60,
         constructing_unit_Datapath_Middle_registers0_h_4_n59,
         constructing_unit_Datapath_Middle_registers0_h_4_n58,
         constructing_unit_Datapath_Middle_registers0_h_4_n57,
         constructing_unit_Datapath_Middle_registers0_h_4_n56,
         constructing_unit_Datapath_Middle_registers0_h_4_n55,
         constructing_unit_Datapath_Middle_registers0_h_4_n54,
         constructing_unit_Datapath_Middle_registers0_h_4_n53,
         constructing_unit_Datapath_Middle_registers0_h_4_n52,
         constructing_unit_Datapath_Middle_registers0_h_4_n51,
         constructing_unit_Datapath_Middle_registers0_h_4_n50,
         constructing_unit_Datapath_Middle_registers0_h_4_n49,
         constructing_unit_Datapath_Middle_registers0_h_4_n48,
         constructing_unit_Datapath_Middle_registers0_h_4_n47,
         constructing_unit_Datapath_Middle_registers0_h_4_n46,
         constructing_unit_Datapath_Middle_registers0_h_4_n45,
         constructing_unit_Datapath_Middle_registers0_h_4_n44,
         constructing_unit_Datapath_Middle_registers0_h_4_n43,
         constructing_unit_Datapath_Middle_registers0_h_4_n42,
         constructing_unit_Datapath_Middle_registers0_h_4_n41,
         constructing_unit_Datapath_Middle_registers0_h_4_n40,
         constructing_unit_Datapath_Middle_registers0_h_4_n39,
         constructing_unit_Datapath_Middle_registers0_h_4_n38,
         constructing_unit_Datapath_Middle_registers0_h_4_n37,
         constructing_unit_Datapath_Middle_registers0_h_4_n36,
         constructing_unit_Datapath_Middle_registers0_h_4_n35,
         constructing_unit_Datapath_Middle_registers0_h_4_n33,
         constructing_unit_Datapath_Middle_registers0_h_5_n67,
         constructing_unit_Datapath_Middle_registers0_h_5_n66,
         constructing_unit_Datapath_Middle_registers0_h_5_n65,
         constructing_unit_Datapath_Middle_registers0_h_5_n64,
         constructing_unit_Datapath_Middle_registers0_h_5_n63,
         constructing_unit_Datapath_Middle_registers0_h_5_n62,
         constructing_unit_Datapath_Middle_registers0_h_5_n61,
         constructing_unit_Datapath_Middle_registers0_h_5_n60,
         constructing_unit_Datapath_Middle_registers0_h_5_n59,
         constructing_unit_Datapath_Middle_registers0_h_5_n58,
         constructing_unit_Datapath_Middle_registers0_h_5_n57,
         constructing_unit_Datapath_Middle_registers0_h_5_n56,
         constructing_unit_Datapath_Middle_registers0_h_5_n55,
         constructing_unit_Datapath_Middle_registers0_h_5_n54,
         constructing_unit_Datapath_Middle_registers0_h_5_n53,
         constructing_unit_Datapath_Middle_registers0_h_5_n52,
         constructing_unit_Datapath_Middle_registers0_h_5_n51,
         constructing_unit_Datapath_Middle_registers0_h_5_n50,
         constructing_unit_Datapath_Middle_registers0_h_5_n49,
         constructing_unit_Datapath_Middle_registers0_h_5_n48,
         constructing_unit_Datapath_Middle_registers0_h_5_n47,
         constructing_unit_Datapath_Middle_registers0_h_5_n46,
         constructing_unit_Datapath_Middle_registers0_h_5_n45,
         constructing_unit_Datapath_Middle_registers0_h_5_n44,
         constructing_unit_Datapath_Middle_registers0_h_5_n43,
         constructing_unit_Datapath_Middle_registers0_h_5_n42,
         constructing_unit_Datapath_Middle_registers0_h_5_n41,
         constructing_unit_Datapath_Middle_registers0_h_5_n40,
         constructing_unit_Datapath_Middle_registers0_h_5_n39,
         constructing_unit_Datapath_Middle_registers0_h_5_n38,
         constructing_unit_Datapath_Middle_registers0_h_5_n37,
         constructing_unit_Datapath_Middle_registers0_h_5_n36,
         constructing_unit_Datapath_Middle_registers0_h_5_n35,
         constructing_unit_Datapath_Middle_registers0_h_5_n33,
         constructing_unit_Datapath_Middle_registers0_h_6_n67,
         constructing_unit_Datapath_Middle_registers0_h_6_n66,
         constructing_unit_Datapath_Middle_registers0_h_6_n65,
         constructing_unit_Datapath_Middle_registers0_h_6_n64,
         constructing_unit_Datapath_Middle_registers0_h_6_n63,
         constructing_unit_Datapath_Middle_registers0_h_6_n62,
         constructing_unit_Datapath_Middle_registers0_h_6_n61,
         constructing_unit_Datapath_Middle_registers0_h_6_n60,
         constructing_unit_Datapath_Middle_registers0_h_6_n59,
         constructing_unit_Datapath_Middle_registers0_h_6_n58,
         constructing_unit_Datapath_Middle_registers0_h_6_n57,
         constructing_unit_Datapath_Middle_registers0_h_6_n56,
         constructing_unit_Datapath_Middle_registers0_h_6_n55,
         constructing_unit_Datapath_Middle_registers0_h_6_n54,
         constructing_unit_Datapath_Middle_registers0_h_6_n53,
         constructing_unit_Datapath_Middle_registers0_h_6_n52,
         constructing_unit_Datapath_Middle_registers0_h_6_n51,
         constructing_unit_Datapath_Middle_registers0_h_6_n50,
         constructing_unit_Datapath_Middle_registers0_h_6_n49,
         constructing_unit_Datapath_Middle_registers0_h_6_n48,
         constructing_unit_Datapath_Middle_registers0_h_6_n47,
         constructing_unit_Datapath_Middle_registers0_h_6_n46,
         constructing_unit_Datapath_Middle_registers0_h_6_n45,
         constructing_unit_Datapath_Middle_registers0_h_6_n44,
         constructing_unit_Datapath_Middle_registers0_h_6_n43,
         constructing_unit_Datapath_Middle_registers0_h_6_n42,
         constructing_unit_Datapath_Middle_registers0_h_6_n41,
         constructing_unit_Datapath_Middle_registers0_h_6_n40,
         constructing_unit_Datapath_Middle_registers0_h_6_n39,
         constructing_unit_Datapath_Middle_registers0_h_6_n38,
         constructing_unit_Datapath_Middle_registers0_h_6_n37,
         constructing_unit_Datapath_Middle_registers0_h_6_n36,
         constructing_unit_Datapath_Middle_registers0_h_6_n35,
         constructing_unit_Datapath_Middle_registers0_h_6_n33,
         constructing_unit_Datapath_Middle_registers0_h_7_n67,
         constructing_unit_Datapath_Middle_registers0_h_7_n66,
         constructing_unit_Datapath_Middle_registers0_h_7_n65,
         constructing_unit_Datapath_Middle_registers0_h_7_n64,
         constructing_unit_Datapath_Middle_registers0_h_7_n63,
         constructing_unit_Datapath_Middle_registers0_h_7_n62,
         constructing_unit_Datapath_Middle_registers0_h_7_n61,
         constructing_unit_Datapath_Middle_registers0_h_7_n60,
         constructing_unit_Datapath_Middle_registers0_h_7_n59,
         constructing_unit_Datapath_Middle_registers0_h_7_n58,
         constructing_unit_Datapath_Middle_registers0_h_7_n57,
         constructing_unit_Datapath_Middle_registers0_h_7_n56,
         constructing_unit_Datapath_Middle_registers0_h_7_n55,
         constructing_unit_Datapath_Middle_registers0_h_7_n54,
         constructing_unit_Datapath_Middle_registers0_h_7_n53,
         constructing_unit_Datapath_Middle_registers0_h_7_n52,
         constructing_unit_Datapath_Middle_registers0_h_7_n51,
         constructing_unit_Datapath_Middle_registers0_h_7_n50,
         constructing_unit_Datapath_Middle_registers0_h_7_n49,
         constructing_unit_Datapath_Middle_registers0_h_7_n48,
         constructing_unit_Datapath_Middle_registers0_h_7_n47,
         constructing_unit_Datapath_Middle_registers0_h_7_n46,
         constructing_unit_Datapath_Middle_registers0_h_7_n45,
         constructing_unit_Datapath_Middle_registers0_h_7_n44,
         constructing_unit_Datapath_Middle_registers0_h_7_n43,
         constructing_unit_Datapath_Middle_registers0_h_7_n42,
         constructing_unit_Datapath_Middle_registers0_h_7_n41,
         constructing_unit_Datapath_Middle_registers0_h_7_n40,
         constructing_unit_Datapath_Middle_registers0_h_7_n39,
         constructing_unit_Datapath_Middle_registers0_h_7_n38,
         constructing_unit_Datapath_Middle_registers0_h_7_n37,
         constructing_unit_Datapath_Middle_registers0_h_7_n36,
         constructing_unit_Datapath_Middle_registers0_h_7_n35,
         constructing_unit_Datapath_Middle_registers0_h_7_n33,
         constructing_unit_Datapath_Middle_registers0_h_8_n67,
         constructing_unit_Datapath_Middle_registers0_h_8_n66,
         constructing_unit_Datapath_Middle_registers0_h_8_n65,
         constructing_unit_Datapath_Middle_registers0_h_8_n64,
         constructing_unit_Datapath_Middle_registers0_h_8_n63,
         constructing_unit_Datapath_Middle_registers0_h_8_n62,
         constructing_unit_Datapath_Middle_registers0_h_8_n61,
         constructing_unit_Datapath_Middle_registers0_h_8_n60,
         constructing_unit_Datapath_Middle_registers0_h_8_n59,
         constructing_unit_Datapath_Middle_registers0_h_8_n58,
         constructing_unit_Datapath_Middle_registers0_h_8_n57,
         constructing_unit_Datapath_Middle_registers0_h_8_n56,
         constructing_unit_Datapath_Middle_registers0_h_8_n55,
         constructing_unit_Datapath_Middle_registers0_h_8_n54,
         constructing_unit_Datapath_Middle_registers0_h_8_n53,
         constructing_unit_Datapath_Middle_registers0_h_8_n52,
         constructing_unit_Datapath_Middle_registers0_h_8_n51,
         constructing_unit_Datapath_Middle_registers0_h_8_n50,
         constructing_unit_Datapath_Middle_registers0_h_8_n49,
         constructing_unit_Datapath_Middle_registers0_h_8_n48,
         constructing_unit_Datapath_Middle_registers0_h_8_n47,
         constructing_unit_Datapath_Middle_registers0_h_8_n46,
         constructing_unit_Datapath_Middle_registers0_h_8_n45,
         constructing_unit_Datapath_Middle_registers0_h_8_n44,
         constructing_unit_Datapath_Middle_registers0_h_8_n43,
         constructing_unit_Datapath_Middle_registers0_h_8_n42,
         constructing_unit_Datapath_Middle_registers0_h_8_n41,
         constructing_unit_Datapath_Middle_registers0_h_8_n40,
         constructing_unit_Datapath_Middle_registers0_h_8_n39,
         constructing_unit_Datapath_Middle_registers0_h_8_n38,
         constructing_unit_Datapath_Middle_registers0_h_8_n37,
         constructing_unit_Datapath_Middle_registers0_h_8_n36,
         constructing_unit_Datapath_Middle_registers0_h_8_n35,
         constructing_unit_Datapath_Middle_registers0_h_8_n33,
         constructing_unit_Datapath_Middle_registers0_h_9_n67,
         constructing_unit_Datapath_Middle_registers0_h_9_n66,
         constructing_unit_Datapath_Middle_registers0_h_9_n65,
         constructing_unit_Datapath_Middle_registers0_h_9_n64,
         constructing_unit_Datapath_Middle_registers0_h_9_n63,
         constructing_unit_Datapath_Middle_registers0_h_9_n62,
         constructing_unit_Datapath_Middle_registers0_h_9_n61,
         constructing_unit_Datapath_Middle_registers0_h_9_n60,
         constructing_unit_Datapath_Middle_registers0_h_9_n59,
         constructing_unit_Datapath_Middle_registers0_h_9_n58,
         constructing_unit_Datapath_Middle_registers0_h_9_n57,
         constructing_unit_Datapath_Middle_registers0_h_9_n56,
         constructing_unit_Datapath_Middle_registers0_h_9_n55,
         constructing_unit_Datapath_Middle_registers0_h_9_n54,
         constructing_unit_Datapath_Middle_registers0_h_9_n53,
         constructing_unit_Datapath_Middle_registers0_h_9_n52,
         constructing_unit_Datapath_Middle_registers0_h_9_n51,
         constructing_unit_Datapath_Middle_registers0_h_9_n50,
         constructing_unit_Datapath_Middle_registers0_h_9_n49,
         constructing_unit_Datapath_Middle_registers0_h_9_n48,
         constructing_unit_Datapath_Middle_registers0_h_9_n47,
         constructing_unit_Datapath_Middle_registers0_h_9_n46,
         constructing_unit_Datapath_Middle_registers0_h_9_n45,
         constructing_unit_Datapath_Middle_registers0_h_9_n44,
         constructing_unit_Datapath_Middle_registers0_h_9_n43,
         constructing_unit_Datapath_Middle_registers0_h_9_n42,
         constructing_unit_Datapath_Middle_registers0_h_9_n41,
         constructing_unit_Datapath_Middle_registers0_h_9_n40,
         constructing_unit_Datapath_Middle_registers0_h_9_n39,
         constructing_unit_Datapath_Middle_registers0_h_9_n38,
         constructing_unit_Datapath_Middle_registers0_h_9_n37,
         constructing_unit_Datapath_Middle_registers0_h_9_n36,
         constructing_unit_Datapath_Middle_registers0_h_9_n35,
         constructing_unit_Datapath_Middle_registers0_h_9_n33,
         constructing_unit_Datapath_Middle_registers0_h_10_n67,
         constructing_unit_Datapath_Middle_registers0_h_10_n66,
         constructing_unit_Datapath_Middle_registers0_h_10_n65,
         constructing_unit_Datapath_Middle_registers0_h_10_n64,
         constructing_unit_Datapath_Middle_registers0_h_10_n63,
         constructing_unit_Datapath_Middle_registers0_h_10_n62,
         constructing_unit_Datapath_Middle_registers0_h_10_n61,
         constructing_unit_Datapath_Middle_registers0_h_10_n60,
         constructing_unit_Datapath_Middle_registers0_h_10_n59,
         constructing_unit_Datapath_Middle_registers0_h_10_n58,
         constructing_unit_Datapath_Middle_registers0_h_10_n57,
         constructing_unit_Datapath_Middle_registers0_h_10_n56,
         constructing_unit_Datapath_Middle_registers0_h_10_n55,
         constructing_unit_Datapath_Middle_registers0_h_10_n54,
         constructing_unit_Datapath_Middle_registers0_h_10_n53,
         constructing_unit_Datapath_Middle_registers0_h_10_n52,
         constructing_unit_Datapath_Middle_registers0_h_10_n51,
         constructing_unit_Datapath_Middle_registers0_h_10_n50,
         constructing_unit_Datapath_Middle_registers0_h_10_n49,
         constructing_unit_Datapath_Middle_registers0_h_10_n48,
         constructing_unit_Datapath_Middle_registers0_h_10_n47,
         constructing_unit_Datapath_Middle_registers0_h_10_n46,
         constructing_unit_Datapath_Middle_registers0_h_10_n45,
         constructing_unit_Datapath_Middle_registers0_h_10_n44,
         constructing_unit_Datapath_Middle_registers0_h_10_n43,
         constructing_unit_Datapath_Middle_registers0_h_10_n42,
         constructing_unit_Datapath_Middle_registers0_h_10_n41,
         constructing_unit_Datapath_Middle_registers0_h_10_n40,
         constructing_unit_Datapath_Middle_registers0_h_10_n39,
         constructing_unit_Datapath_Middle_registers0_h_10_n38,
         constructing_unit_Datapath_Middle_registers0_h_10_n37,
         constructing_unit_Datapath_Middle_registers0_h_10_n36,
         constructing_unit_Datapath_Middle_registers0_h_10_n35,
         constructing_unit_Datapath_Middle_registers0_h_10_n33,
         constructing_unit_Datapath_Middle_registers0_h_11_n67,
         constructing_unit_Datapath_Middle_registers0_h_11_n66,
         constructing_unit_Datapath_Middle_registers0_h_11_n65,
         constructing_unit_Datapath_Middle_registers0_h_11_n64,
         constructing_unit_Datapath_Middle_registers0_h_11_n63,
         constructing_unit_Datapath_Middle_registers0_h_11_n62,
         constructing_unit_Datapath_Middle_registers0_h_11_n61,
         constructing_unit_Datapath_Middle_registers0_h_11_n60,
         constructing_unit_Datapath_Middle_registers0_h_11_n59,
         constructing_unit_Datapath_Middle_registers0_h_11_n58,
         constructing_unit_Datapath_Middle_registers0_h_11_n57,
         constructing_unit_Datapath_Middle_registers0_h_11_n56,
         constructing_unit_Datapath_Middle_registers0_h_11_n55,
         constructing_unit_Datapath_Middle_registers0_h_11_n54,
         constructing_unit_Datapath_Middle_registers0_h_11_n53,
         constructing_unit_Datapath_Middle_registers0_h_11_n52,
         constructing_unit_Datapath_Middle_registers0_h_11_n51,
         constructing_unit_Datapath_Middle_registers0_h_11_n50,
         constructing_unit_Datapath_Middle_registers0_h_11_n49,
         constructing_unit_Datapath_Middle_registers0_h_11_n48,
         constructing_unit_Datapath_Middle_registers0_h_11_n47,
         constructing_unit_Datapath_Middle_registers0_h_11_n46,
         constructing_unit_Datapath_Middle_registers0_h_11_n45,
         constructing_unit_Datapath_Middle_registers0_h_11_n44,
         constructing_unit_Datapath_Middle_registers0_h_11_n43,
         constructing_unit_Datapath_Middle_registers0_h_11_n42,
         constructing_unit_Datapath_Middle_registers0_h_11_n41,
         constructing_unit_Datapath_Middle_registers0_h_11_n40,
         constructing_unit_Datapath_Middle_registers0_h_11_n39,
         constructing_unit_Datapath_Middle_registers0_h_11_n38,
         constructing_unit_Datapath_Middle_registers0_h_11_n37,
         constructing_unit_Datapath_Middle_registers0_h_11_n36,
         constructing_unit_Datapath_Middle_registers0_h_11_n35,
         constructing_unit_Datapath_Middle_registers0_h_11_n33,
         constructing_unit_Datapath_Middle_registers0_h_12_n67,
         constructing_unit_Datapath_Middle_registers0_h_12_n66,
         constructing_unit_Datapath_Middle_registers0_h_12_n65,
         constructing_unit_Datapath_Middle_registers0_h_12_n64,
         constructing_unit_Datapath_Middle_registers0_h_12_n63,
         constructing_unit_Datapath_Middle_registers0_h_12_n62,
         constructing_unit_Datapath_Middle_registers0_h_12_n61,
         constructing_unit_Datapath_Middle_registers0_h_12_n60,
         constructing_unit_Datapath_Middle_registers0_h_12_n59,
         constructing_unit_Datapath_Middle_registers0_h_12_n58,
         constructing_unit_Datapath_Middle_registers0_h_12_n57,
         constructing_unit_Datapath_Middle_registers0_h_12_n56,
         constructing_unit_Datapath_Middle_registers0_h_12_n55,
         constructing_unit_Datapath_Middle_registers0_h_12_n54,
         constructing_unit_Datapath_Middle_registers0_h_12_n53,
         constructing_unit_Datapath_Middle_registers0_h_12_n52,
         constructing_unit_Datapath_Middle_registers0_h_12_n51,
         constructing_unit_Datapath_Middle_registers0_h_12_n50,
         constructing_unit_Datapath_Middle_registers0_h_12_n49,
         constructing_unit_Datapath_Middle_registers0_h_12_n48,
         constructing_unit_Datapath_Middle_registers0_h_12_n47,
         constructing_unit_Datapath_Middle_registers0_h_12_n46,
         constructing_unit_Datapath_Middle_registers0_h_12_n45,
         constructing_unit_Datapath_Middle_registers0_h_12_n44,
         constructing_unit_Datapath_Middle_registers0_h_12_n43,
         constructing_unit_Datapath_Middle_registers0_h_12_n42,
         constructing_unit_Datapath_Middle_registers0_h_12_n41,
         constructing_unit_Datapath_Middle_registers0_h_12_n40,
         constructing_unit_Datapath_Middle_registers0_h_12_n39,
         constructing_unit_Datapath_Middle_registers0_h_12_n38,
         constructing_unit_Datapath_Middle_registers0_h_12_n37,
         constructing_unit_Datapath_Middle_registers0_h_12_n36,
         constructing_unit_Datapath_Middle_registers0_h_12_n35,
         constructing_unit_Datapath_Middle_registers0_h_12_n33,
         constructing_unit_Datapath_Middle_registers0_h_13_n67,
         constructing_unit_Datapath_Middle_registers0_h_13_n66,
         constructing_unit_Datapath_Middle_registers0_h_13_n65,
         constructing_unit_Datapath_Middle_registers0_h_13_n64,
         constructing_unit_Datapath_Middle_registers0_h_13_n63,
         constructing_unit_Datapath_Middle_registers0_h_13_n62,
         constructing_unit_Datapath_Middle_registers0_h_13_n61,
         constructing_unit_Datapath_Middle_registers0_h_13_n60,
         constructing_unit_Datapath_Middle_registers0_h_13_n59,
         constructing_unit_Datapath_Middle_registers0_h_13_n58,
         constructing_unit_Datapath_Middle_registers0_h_13_n57,
         constructing_unit_Datapath_Middle_registers0_h_13_n56,
         constructing_unit_Datapath_Middle_registers0_h_13_n55,
         constructing_unit_Datapath_Middle_registers0_h_13_n54,
         constructing_unit_Datapath_Middle_registers0_h_13_n53,
         constructing_unit_Datapath_Middle_registers0_h_13_n52,
         constructing_unit_Datapath_Middle_registers0_h_13_n51,
         constructing_unit_Datapath_Middle_registers0_h_13_n50,
         constructing_unit_Datapath_Middle_registers0_h_13_n49,
         constructing_unit_Datapath_Middle_registers0_h_13_n48,
         constructing_unit_Datapath_Middle_registers0_h_13_n47,
         constructing_unit_Datapath_Middle_registers0_h_13_n46,
         constructing_unit_Datapath_Middle_registers0_h_13_n45,
         constructing_unit_Datapath_Middle_registers0_h_13_n44,
         constructing_unit_Datapath_Middle_registers0_h_13_n43,
         constructing_unit_Datapath_Middle_registers0_h_13_n42,
         constructing_unit_Datapath_Middle_registers0_h_13_n41,
         constructing_unit_Datapath_Middle_registers0_h_13_n40,
         constructing_unit_Datapath_Middle_registers0_h_13_n39,
         constructing_unit_Datapath_Middle_registers0_h_13_n38,
         constructing_unit_Datapath_Middle_registers0_h_13_n37,
         constructing_unit_Datapath_Middle_registers0_h_13_n36,
         constructing_unit_Datapath_Middle_registers0_h_13_n35,
         constructing_unit_Datapath_Middle_registers0_h_13_n33,
         constructing_unit_Datapath_Middle_registers1_3_n67,
         constructing_unit_Datapath_Middle_registers1_3_n66,
         constructing_unit_Datapath_Middle_registers1_3_n65,
         constructing_unit_Datapath_Middle_registers1_3_n64,
         constructing_unit_Datapath_Middle_registers1_3_n63,
         constructing_unit_Datapath_Middle_registers1_3_n62,
         constructing_unit_Datapath_Middle_registers1_3_n61,
         constructing_unit_Datapath_Middle_registers1_3_n60,
         constructing_unit_Datapath_Middle_registers1_3_n59,
         constructing_unit_Datapath_Middle_registers1_3_n58,
         constructing_unit_Datapath_Middle_registers1_3_n57,
         constructing_unit_Datapath_Middle_registers1_3_n56,
         constructing_unit_Datapath_Middle_registers1_3_n55,
         constructing_unit_Datapath_Middle_registers1_3_n54,
         constructing_unit_Datapath_Middle_registers1_3_n53,
         constructing_unit_Datapath_Middle_registers1_3_n52,
         constructing_unit_Datapath_Middle_registers1_3_n51,
         constructing_unit_Datapath_Middle_registers1_3_n50,
         constructing_unit_Datapath_Middle_registers1_3_n49,
         constructing_unit_Datapath_Middle_registers1_3_n48,
         constructing_unit_Datapath_Middle_registers1_3_n47,
         constructing_unit_Datapath_Middle_registers1_3_n46,
         constructing_unit_Datapath_Middle_registers1_3_n45,
         constructing_unit_Datapath_Middle_registers1_3_n44,
         constructing_unit_Datapath_Middle_registers1_3_n43,
         constructing_unit_Datapath_Middle_registers1_3_n42,
         constructing_unit_Datapath_Middle_registers1_3_n41,
         constructing_unit_Datapath_Middle_registers1_3_n40,
         constructing_unit_Datapath_Middle_registers1_3_n39,
         constructing_unit_Datapath_Middle_registers1_3_n38,
         constructing_unit_Datapath_Middle_registers1_3_n37,
         constructing_unit_Datapath_Middle_registers1_3_n36,
         constructing_unit_Datapath_Middle_registers1_3_n35,
         constructing_unit_Datapath_Middle_registers1_3_n33,
         constructing_unit_Datapath_Middle_registers1_4_n67,
         constructing_unit_Datapath_Middle_registers1_4_n66,
         constructing_unit_Datapath_Middle_registers1_4_n65,
         constructing_unit_Datapath_Middle_registers1_4_n64,
         constructing_unit_Datapath_Middle_registers1_4_n63,
         constructing_unit_Datapath_Middle_registers1_4_n62,
         constructing_unit_Datapath_Middle_registers1_4_n61,
         constructing_unit_Datapath_Middle_registers1_4_n60,
         constructing_unit_Datapath_Middle_registers1_4_n59,
         constructing_unit_Datapath_Middle_registers1_4_n58,
         constructing_unit_Datapath_Middle_registers1_4_n57,
         constructing_unit_Datapath_Middle_registers1_4_n56,
         constructing_unit_Datapath_Middle_registers1_4_n55,
         constructing_unit_Datapath_Middle_registers1_4_n54,
         constructing_unit_Datapath_Middle_registers1_4_n53,
         constructing_unit_Datapath_Middle_registers1_4_n52,
         constructing_unit_Datapath_Middle_registers1_4_n51,
         constructing_unit_Datapath_Middle_registers1_4_n50,
         constructing_unit_Datapath_Middle_registers1_4_n49,
         constructing_unit_Datapath_Middle_registers1_4_n48,
         constructing_unit_Datapath_Middle_registers1_4_n47,
         constructing_unit_Datapath_Middle_registers1_4_n46,
         constructing_unit_Datapath_Middle_registers1_4_n45,
         constructing_unit_Datapath_Middle_registers1_4_n44,
         constructing_unit_Datapath_Middle_registers1_4_n43,
         constructing_unit_Datapath_Middle_registers1_4_n42,
         constructing_unit_Datapath_Middle_registers1_4_n41,
         constructing_unit_Datapath_Middle_registers1_4_n40,
         constructing_unit_Datapath_Middle_registers1_4_n39,
         constructing_unit_Datapath_Middle_registers1_4_n38,
         constructing_unit_Datapath_Middle_registers1_4_n37,
         constructing_unit_Datapath_Middle_registers1_4_n36,
         constructing_unit_Datapath_Middle_registers1_4_n35,
         constructing_unit_Datapath_Middle_registers1_4_n33,
         constructing_unit_Datapath_Middle_registers1_5_n67,
         constructing_unit_Datapath_Middle_registers1_5_n66,
         constructing_unit_Datapath_Middle_registers1_5_n65,
         constructing_unit_Datapath_Middle_registers1_5_n64,
         constructing_unit_Datapath_Middle_registers1_5_n63,
         constructing_unit_Datapath_Middle_registers1_5_n62,
         constructing_unit_Datapath_Middle_registers1_5_n61,
         constructing_unit_Datapath_Middle_registers1_5_n60,
         constructing_unit_Datapath_Middle_registers1_5_n59,
         constructing_unit_Datapath_Middle_registers1_5_n58,
         constructing_unit_Datapath_Middle_registers1_5_n57,
         constructing_unit_Datapath_Middle_registers1_5_n56,
         constructing_unit_Datapath_Middle_registers1_5_n55,
         constructing_unit_Datapath_Middle_registers1_5_n54,
         constructing_unit_Datapath_Middle_registers1_5_n53,
         constructing_unit_Datapath_Middle_registers1_5_n52,
         constructing_unit_Datapath_Middle_registers1_5_n51,
         constructing_unit_Datapath_Middle_registers1_5_n50,
         constructing_unit_Datapath_Middle_registers1_5_n49,
         constructing_unit_Datapath_Middle_registers1_5_n48,
         constructing_unit_Datapath_Middle_registers1_5_n47,
         constructing_unit_Datapath_Middle_registers1_5_n46,
         constructing_unit_Datapath_Middle_registers1_5_n45,
         constructing_unit_Datapath_Middle_registers1_5_n44,
         constructing_unit_Datapath_Middle_registers1_5_n43,
         constructing_unit_Datapath_Middle_registers1_5_n42,
         constructing_unit_Datapath_Middle_registers1_5_n41,
         constructing_unit_Datapath_Middle_registers1_5_n40,
         constructing_unit_Datapath_Middle_registers1_5_n39,
         constructing_unit_Datapath_Middle_registers1_5_n38,
         constructing_unit_Datapath_Middle_registers1_5_n37,
         constructing_unit_Datapath_Middle_registers1_5_n36,
         constructing_unit_Datapath_Middle_registers1_5_n35,
         constructing_unit_Datapath_Middle_registers1_5_n33,
         constructing_unit_Datapath_Middle_registers1_6_n67,
         constructing_unit_Datapath_Middle_registers1_6_n66,
         constructing_unit_Datapath_Middle_registers1_6_n65,
         constructing_unit_Datapath_Middle_registers1_6_n64,
         constructing_unit_Datapath_Middle_registers1_6_n63,
         constructing_unit_Datapath_Middle_registers1_6_n62,
         constructing_unit_Datapath_Middle_registers1_6_n61,
         constructing_unit_Datapath_Middle_registers1_6_n60,
         constructing_unit_Datapath_Middle_registers1_6_n59,
         constructing_unit_Datapath_Middle_registers1_6_n58,
         constructing_unit_Datapath_Middle_registers1_6_n57,
         constructing_unit_Datapath_Middle_registers1_6_n56,
         constructing_unit_Datapath_Middle_registers1_6_n55,
         constructing_unit_Datapath_Middle_registers1_6_n54,
         constructing_unit_Datapath_Middle_registers1_6_n53,
         constructing_unit_Datapath_Middle_registers1_6_n52,
         constructing_unit_Datapath_Middle_registers1_6_n51,
         constructing_unit_Datapath_Middle_registers1_6_n50,
         constructing_unit_Datapath_Middle_registers1_6_n49,
         constructing_unit_Datapath_Middle_registers1_6_n48,
         constructing_unit_Datapath_Middle_registers1_6_n47,
         constructing_unit_Datapath_Middle_registers1_6_n46,
         constructing_unit_Datapath_Middle_registers1_6_n45,
         constructing_unit_Datapath_Middle_registers1_6_n44,
         constructing_unit_Datapath_Middle_registers1_6_n43,
         constructing_unit_Datapath_Middle_registers1_6_n42,
         constructing_unit_Datapath_Middle_registers1_6_n41,
         constructing_unit_Datapath_Middle_registers1_6_n40,
         constructing_unit_Datapath_Middle_registers1_6_n39,
         constructing_unit_Datapath_Middle_registers1_6_n38,
         constructing_unit_Datapath_Middle_registers1_6_n37,
         constructing_unit_Datapath_Middle_registers1_6_n36,
         constructing_unit_Datapath_Middle_registers1_6_n35,
         constructing_unit_Datapath_Middle_registers1_6_n33,
         constructing_unit_Datapath_Middle_registers1_7_n67,
         constructing_unit_Datapath_Middle_registers1_7_n66,
         constructing_unit_Datapath_Middle_registers1_7_n65,
         constructing_unit_Datapath_Middle_registers1_7_n64,
         constructing_unit_Datapath_Middle_registers1_7_n63,
         constructing_unit_Datapath_Middle_registers1_7_n62,
         constructing_unit_Datapath_Middle_registers1_7_n61,
         constructing_unit_Datapath_Middle_registers1_7_n60,
         constructing_unit_Datapath_Middle_registers1_7_n59,
         constructing_unit_Datapath_Middle_registers1_7_n58,
         constructing_unit_Datapath_Middle_registers1_7_n57,
         constructing_unit_Datapath_Middle_registers1_7_n56,
         constructing_unit_Datapath_Middle_registers1_7_n55,
         constructing_unit_Datapath_Middle_registers1_7_n54,
         constructing_unit_Datapath_Middle_registers1_7_n53,
         constructing_unit_Datapath_Middle_registers1_7_n52,
         constructing_unit_Datapath_Middle_registers1_7_n51,
         constructing_unit_Datapath_Middle_registers1_7_n50,
         constructing_unit_Datapath_Middle_registers1_7_n49,
         constructing_unit_Datapath_Middle_registers1_7_n48,
         constructing_unit_Datapath_Middle_registers1_7_n47,
         constructing_unit_Datapath_Middle_registers1_7_n46,
         constructing_unit_Datapath_Middle_registers1_7_n45,
         constructing_unit_Datapath_Middle_registers1_7_n44,
         constructing_unit_Datapath_Middle_registers1_7_n43,
         constructing_unit_Datapath_Middle_registers1_7_n42,
         constructing_unit_Datapath_Middle_registers1_7_n41,
         constructing_unit_Datapath_Middle_registers1_7_n40,
         constructing_unit_Datapath_Middle_registers1_7_n39,
         constructing_unit_Datapath_Middle_registers1_7_n38,
         constructing_unit_Datapath_Middle_registers1_7_n37,
         constructing_unit_Datapath_Middle_registers1_7_n36,
         constructing_unit_Datapath_Middle_registers1_7_n35,
         constructing_unit_Datapath_Middle_registers1_7_n33,
         constructing_unit_Datapath_Middle_registers1_8_n67,
         constructing_unit_Datapath_Middle_registers1_8_n66,
         constructing_unit_Datapath_Middle_registers1_8_n65,
         constructing_unit_Datapath_Middle_registers1_8_n64,
         constructing_unit_Datapath_Middle_registers1_8_n63,
         constructing_unit_Datapath_Middle_registers1_8_n62,
         constructing_unit_Datapath_Middle_registers1_8_n61,
         constructing_unit_Datapath_Middle_registers1_8_n60,
         constructing_unit_Datapath_Middle_registers1_8_n59,
         constructing_unit_Datapath_Middle_registers1_8_n58,
         constructing_unit_Datapath_Middle_registers1_8_n57,
         constructing_unit_Datapath_Middle_registers1_8_n56,
         constructing_unit_Datapath_Middle_registers1_8_n55,
         constructing_unit_Datapath_Middle_registers1_8_n54,
         constructing_unit_Datapath_Middle_registers1_8_n53,
         constructing_unit_Datapath_Middle_registers1_8_n52,
         constructing_unit_Datapath_Middle_registers1_8_n51,
         constructing_unit_Datapath_Middle_registers1_8_n50,
         constructing_unit_Datapath_Middle_registers1_8_n49,
         constructing_unit_Datapath_Middle_registers1_8_n48,
         constructing_unit_Datapath_Middle_registers1_8_n47,
         constructing_unit_Datapath_Middle_registers1_8_n46,
         constructing_unit_Datapath_Middle_registers1_8_n45,
         constructing_unit_Datapath_Middle_registers1_8_n44,
         constructing_unit_Datapath_Middle_registers1_8_n43,
         constructing_unit_Datapath_Middle_registers1_8_n42,
         constructing_unit_Datapath_Middle_registers1_8_n41,
         constructing_unit_Datapath_Middle_registers1_8_n40,
         constructing_unit_Datapath_Middle_registers1_8_n39,
         constructing_unit_Datapath_Middle_registers1_8_n38,
         constructing_unit_Datapath_Middle_registers1_8_n37,
         constructing_unit_Datapath_Middle_registers1_8_n36,
         constructing_unit_Datapath_Middle_registers1_8_n35,
         constructing_unit_Datapath_Middle_registers1_8_n33,
         constructing_unit_Datapath_Middle_registers1_9_n67,
         constructing_unit_Datapath_Middle_registers1_9_n66,
         constructing_unit_Datapath_Middle_registers1_9_n65,
         constructing_unit_Datapath_Middle_registers1_9_n64,
         constructing_unit_Datapath_Middle_registers1_9_n63,
         constructing_unit_Datapath_Middle_registers1_9_n62,
         constructing_unit_Datapath_Middle_registers1_9_n61,
         constructing_unit_Datapath_Middle_registers1_9_n60,
         constructing_unit_Datapath_Middle_registers1_9_n59,
         constructing_unit_Datapath_Middle_registers1_9_n58,
         constructing_unit_Datapath_Middle_registers1_9_n57,
         constructing_unit_Datapath_Middle_registers1_9_n56,
         constructing_unit_Datapath_Middle_registers1_9_n55,
         constructing_unit_Datapath_Middle_registers1_9_n54,
         constructing_unit_Datapath_Middle_registers1_9_n53,
         constructing_unit_Datapath_Middle_registers1_9_n52,
         constructing_unit_Datapath_Middle_registers1_9_n51,
         constructing_unit_Datapath_Middle_registers1_9_n50,
         constructing_unit_Datapath_Middle_registers1_9_n49,
         constructing_unit_Datapath_Middle_registers1_9_n48,
         constructing_unit_Datapath_Middle_registers1_9_n47,
         constructing_unit_Datapath_Middle_registers1_9_n46,
         constructing_unit_Datapath_Middle_registers1_9_n45,
         constructing_unit_Datapath_Middle_registers1_9_n44,
         constructing_unit_Datapath_Middle_registers1_9_n43,
         constructing_unit_Datapath_Middle_registers1_9_n42,
         constructing_unit_Datapath_Middle_registers1_9_n41,
         constructing_unit_Datapath_Middle_registers1_9_n40,
         constructing_unit_Datapath_Middle_registers1_9_n39,
         constructing_unit_Datapath_Middle_registers1_9_n38,
         constructing_unit_Datapath_Middle_registers1_9_n37,
         constructing_unit_Datapath_Middle_registers1_9_n36,
         constructing_unit_Datapath_Middle_registers1_9_n35,
         constructing_unit_Datapath_Middle_registers1_9_n33,
         constructing_unit_Datapath_Middle_registers1_10_n67,
         constructing_unit_Datapath_Middle_registers1_10_n66,
         constructing_unit_Datapath_Middle_registers1_10_n65,
         constructing_unit_Datapath_Middle_registers1_10_n64,
         constructing_unit_Datapath_Middle_registers1_10_n63,
         constructing_unit_Datapath_Middle_registers1_10_n62,
         constructing_unit_Datapath_Middle_registers1_10_n61,
         constructing_unit_Datapath_Middle_registers1_10_n60,
         constructing_unit_Datapath_Middle_registers1_10_n59,
         constructing_unit_Datapath_Middle_registers1_10_n58,
         constructing_unit_Datapath_Middle_registers1_10_n57,
         constructing_unit_Datapath_Middle_registers1_10_n56,
         constructing_unit_Datapath_Middle_registers1_10_n55,
         constructing_unit_Datapath_Middle_registers1_10_n54,
         constructing_unit_Datapath_Middle_registers1_10_n53,
         constructing_unit_Datapath_Middle_registers1_10_n52,
         constructing_unit_Datapath_Middle_registers1_10_n51,
         constructing_unit_Datapath_Middle_registers1_10_n50,
         constructing_unit_Datapath_Middle_registers1_10_n49,
         constructing_unit_Datapath_Middle_registers1_10_n48,
         constructing_unit_Datapath_Middle_registers1_10_n47,
         constructing_unit_Datapath_Middle_registers1_10_n46,
         constructing_unit_Datapath_Middle_registers1_10_n45,
         constructing_unit_Datapath_Middle_registers1_10_n44,
         constructing_unit_Datapath_Middle_registers1_10_n43,
         constructing_unit_Datapath_Middle_registers1_10_n42,
         constructing_unit_Datapath_Middle_registers1_10_n41,
         constructing_unit_Datapath_Middle_registers1_10_n40,
         constructing_unit_Datapath_Middle_registers1_10_n39,
         constructing_unit_Datapath_Middle_registers1_10_n38,
         constructing_unit_Datapath_Middle_registers1_10_n37,
         constructing_unit_Datapath_Middle_registers1_10_n36,
         constructing_unit_Datapath_Middle_registers1_10_n35,
         constructing_unit_Datapath_Middle_registers1_10_n33,
         constructing_unit_Datapath_Middle_registers1_11_n67,
         constructing_unit_Datapath_Middle_registers1_11_n66,
         constructing_unit_Datapath_Middle_registers1_11_n65,
         constructing_unit_Datapath_Middle_registers1_11_n64,
         constructing_unit_Datapath_Middle_registers1_11_n63,
         constructing_unit_Datapath_Middle_registers1_11_n62,
         constructing_unit_Datapath_Middle_registers1_11_n61,
         constructing_unit_Datapath_Middle_registers1_11_n60,
         constructing_unit_Datapath_Middle_registers1_11_n59,
         constructing_unit_Datapath_Middle_registers1_11_n58,
         constructing_unit_Datapath_Middle_registers1_11_n57,
         constructing_unit_Datapath_Middle_registers1_11_n56,
         constructing_unit_Datapath_Middle_registers1_11_n55,
         constructing_unit_Datapath_Middle_registers1_11_n54,
         constructing_unit_Datapath_Middle_registers1_11_n53,
         constructing_unit_Datapath_Middle_registers1_11_n52,
         constructing_unit_Datapath_Middle_registers1_11_n51,
         constructing_unit_Datapath_Middle_registers1_11_n50,
         constructing_unit_Datapath_Middle_registers1_11_n49,
         constructing_unit_Datapath_Middle_registers1_11_n48,
         constructing_unit_Datapath_Middle_registers1_11_n47,
         constructing_unit_Datapath_Middle_registers1_11_n46,
         constructing_unit_Datapath_Middle_registers1_11_n45,
         constructing_unit_Datapath_Middle_registers1_11_n44,
         constructing_unit_Datapath_Middle_registers1_11_n43,
         constructing_unit_Datapath_Middle_registers1_11_n42,
         constructing_unit_Datapath_Middle_registers1_11_n41,
         constructing_unit_Datapath_Middle_registers1_11_n40,
         constructing_unit_Datapath_Middle_registers1_11_n39,
         constructing_unit_Datapath_Middle_registers1_11_n38,
         constructing_unit_Datapath_Middle_registers1_11_n37,
         constructing_unit_Datapath_Middle_registers1_11_n36,
         constructing_unit_Datapath_Middle_registers1_11_n35,
         constructing_unit_Datapath_Middle_registers1_11_n33,
         constructing_unit_Datapath_Middle_registers1_12_n67,
         constructing_unit_Datapath_Middle_registers1_12_n66,
         constructing_unit_Datapath_Middle_registers1_12_n65,
         constructing_unit_Datapath_Middle_registers1_12_n64,
         constructing_unit_Datapath_Middle_registers1_12_n63,
         constructing_unit_Datapath_Middle_registers1_12_n62,
         constructing_unit_Datapath_Middle_registers1_12_n61,
         constructing_unit_Datapath_Middle_registers1_12_n60,
         constructing_unit_Datapath_Middle_registers1_12_n59,
         constructing_unit_Datapath_Middle_registers1_12_n58,
         constructing_unit_Datapath_Middle_registers1_12_n57,
         constructing_unit_Datapath_Middle_registers1_12_n56,
         constructing_unit_Datapath_Middle_registers1_12_n55,
         constructing_unit_Datapath_Middle_registers1_12_n54,
         constructing_unit_Datapath_Middle_registers1_12_n53,
         constructing_unit_Datapath_Middle_registers1_12_n52,
         constructing_unit_Datapath_Middle_registers1_12_n51,
         constructing_unit_Datapath_Middle_registers1_12_n50,
         constructing_unit_Datapath_Middle_registers1_12_n49,
         constructing_unit_Datapath_Middle_registers1_12_n48,
         constructing_unit_Datapath_Middle_registers1_12_n47,
         constructing_unit_Datapath_Middle_registers1_12_n46,
         constructing_unit_Datapath_Middle_registers1_12_n45,
         constructing_unit_Datapath_Middle_registers1_12_n44,
         constructing_unit_Datapath_Middle_registers1_12_n43,
         constructing_unit_Datapath_Middle_registers1_12_n42,
         constructing_unit_Datapath_Middle_registers1_12_n41,
         constructing_unit_Datapath_Middle_registers1_12_n40,
         constructing_unit_Datapath_Middle_registers1_12_n39,
         constructing_unit_Datapath_Middle_registers1_12_n38,
         constructing_unit_Datapath_Middle_registers1_12_n37,
         constructing_unit_Datapath_Middle_registers1_12_n36,
         constructing_unit_Datapath_Middle_registers1_12_n35,
         constructing_unit_Datapath_Middle_registers1_12_n33,
         constructing_unit_Datapath_Middle_registers1_13_n67,
         constructing_unit_Datapath_Middle_registers1_13_n66,
         constructing_unit_Datapath_Middle_registers1_13_n65,
         constructing_unit_Datapath_Middle_registers1_13_n64,
         constructing_unit_Datapath_Middle_registers1_13_n63,
         constructing_unit_Datapath_Middle_registers1_13_n62,
         constructing_unit_Datapath_Middle_registers1_13_n61,
         constructing_unit_Datapath_Middle_registers1_13_n60,
         constructing_unit_Datapath_Middle_registers1_13_n59,
         constructing_unit_Datapath_Middle_registers1_13_n58,
         constructing_unit_Datapath_Middle_registers1_13_n57,
         constructing_unit_Datapath_Middle_registers1_13_n56,
         constructing_unit_Datapath_Middle_registers1_13_n55,
         constructing_unit_Datapath_Middle_registers1_13_n54,
         constructing_unit_Datapath_Middle_registers1_13_n53,
         constructing_unit_Datapath_Middle_registers1_13_n52,
         constructing_unit_Datapath_Middle_registers1_13_n51,
         constructing_unit_Datapath_Middle_registers1_13_n50,
         constructing_unit_Datapath_Middle_registers1_13_n49,
         constructing_unit_Datapath_Middle_registers1_13_n48,
         constructing_unit_Datapath_Middle_registers1_13_n47,
         constructing_unit_Datapath_Middle_registers1_13_n46,
         constructing_unit_Datapath_Middle_registers1_13_n45,
         constructing_unit_Datapath_Middle_registers1_13_n44,
         constructing_unit_Datapath_Middle_registers1_13_n43,
         constructing_unit_Datapath_Middle_registers1_13_n42,
         constructing_unit_Datapath_Middle_registers1_13_n41,
         constructing_unit_Datapath_Middle_registers1_13_n40,
         constructing_unit_Datapath_Middle_registers1_13_n39,
         constructing_unit_Datapath_Middle_registers1_13_n38,
         constructing_unit_Datapath_Middle_registers1_13_n37,
         constructing_unit_Datapath_Middle_registers1_13_n36,
         constructing_unit_Datapath_Middle_registers1_13_n35,
         constructing_unit_Datapath_Middle_registers1_13_n33,
         constructing_unit_Datapath_Middle_registers2_3_n67,
         constructing_unit_Datapath_Middle_registers2_3_n66,
         constructing_unit_Datapath_Middle_registers2_3_n65,
         constructing_unit_Datapath_Middle_registers2_3_n64,
         constructing_unit_Datapath_Middle_registers2_3_n63,
         constructing_unit_Datapath_Middle_registers2_3_n62,
         constructing_unit_Datapath_Middle_registers2_3_n61,
         constructing_unit_Datapath_Middle_registers2_3_n60,
         constructing_unit_Datapath_Middle_registers2_3_n59,
         constructing_unit_Datapath_Middle_registers2_3_n58,
         constructing_unit_Datapath_Middle_registers2_3_n57,
         constructing_unit_Datapath_Middle_registers2_3_n56,
         constructing_unit_Datapath_Middle_registers2_3_n55,
         constructing_unit_Datapath_Middle_registers2_3_n54,
         constructing_unit_Datapath_Middle_registers2_3_n53,
         constructing_unit_Datapath_Middle_registers2_3_n52,
         constructing_unit_Datapath_Middle_registers2_3_n51,
         constructing_unit_Datapath_Middle_registers2_3_n50,
         constructing_unit_Datapath_Middle_registers2_3_n49,
         constructing_unit_Datapath_Middle_registers2_3_n48,
         constructing_unit_Datapath_Middle_registers2_3_n47,
         constructing_unit_Datapath_Middle_registers2_3_n46,
         constructing_unit_Datapath_Middle_registers2_3_n45,
         constructing_unit_Datapath_Middle_registers2_3_n44,
         constructing_unit_Datapath_Middle_registers2_3_n43,
         constructing_unit_Datapath_Middle_registers2_3_n42,
         constructing_unit_Datapath_Middle_registers2_3_n41,
         constructing_unit_Datapath_Middle_registers2_3_n40,
         constructing_unit_Datapath_Middle_registers2_3_n39,
         constructing_unit_Datapath_Middle_registers2_3_n38,
         constructing_unit_Datapath_Middle_registers2_3_n37,
         constructing_unit_Datapath_Middle_registers2_3_n36,
         constructing_unit_Datapath_Middle_registers2_3_n35,
         constructing_unit_Datapath_Middle_registers2_3_n33,
         constructing_unit_Datapath_Middle_registers2_4_n67,
         constructing_unit_Datapath_Middle_registers2_4_n66,
         constructing_unit_Datapath_Middle_registers2_4_n65,
         constructing_unit_Datapath_Middle_registers2_4_n64,
         constructing_unit_Datapath_Middle_registers2_4_n63,
         constructing_unit_Datapath_Middle_registers2_4_n62,
         constructing_unit_Datapath_Middle_registers2_4_n61,
         constructing_unit_Datapath_Middle_registers2_4_n60,
         constructing_unit_Datapath_Middle_registers2_4_n59,
         constructing_unit_Datapath_Middle_registers2_4_n58,
         constructing_unit_Datapath_Middle_registers2_4_n57,
         constructing_unit_Datapath_Middle_registers2_4_n56,
         constructing_unit_Datapath_Middle_registers2_4_n55,
         constructing_unit_Datapath_Middle_registers2_4_n54,
         constructing_unit_Datapath_Middle_registers2_4_n53,
         constructing_unit_Datapath_Middle_registers2_4_n52,
         constructing_unit_Datapath_Middle_registers2_4_n51,
         constructing_unit_Datapath_Middle_registers2_4_n50,
         constructing_unit_Datapath_Middle_registers2_4_n49,
         constructing_unit_Datapath_Middle_registers2_4_n48,
         constructing_unit_Datapath_Middle_registers2_4_n47,
         constructing_unit_Datapath_Middle_registers2_4_n46,
         constructing_unit_Datapath_Middle_registers2_4_n45,
         constructing_unit_Datapath_Middle_registers2_4_n44,
         constructing_unit_Datapath_Middle_registers2_4_n43,
         constructing_unit_Datapath_Middle_registers2_4_n42,
         constructing_unit_Datapath_Middle_registers2_4_n41,
         constructing_unit_Datapath_Middle_registers2_4_n40,
         constructing_unit_Datapath_Middle_registers2_4_n39,
         constructing_unit_Datapath_Middle_registers2_4_n38,
         constructing_unit_Datapath_Middle_registers2_4_n37,
         constructing_unit_Datapath_Middle_registers2_4_n36,
         constructing_unit_Datapath_Middle_registers2_4_n35,
         constructing_unit_Datapath_Middle_registers2_4_n33,
         constructing_unit_Datapath_Middle_registers2_5_n67,
         constructing_unit_Datapath_Middle_registers2_5_n66,
         constructing_unit_Datapath_Middle_registers2_5_n65,
         constructing_unit_Datapath_Middle_registers2_5_n64,
         constructing_unit_Datapath_Middle_registers2_5_n63,
         constructing_unit_Datapath_Middle_registers2_5_n62,
         constructing_unit_Datapath_Middle_registers2_5_n61,
         constructing_unit_Datapath_Middle_registers2_5_n60,
         constructing_unit_Datapath_Middle_registers2_5_n59,
         constructing_unit_Datapath_Middle_registers2_5_n58,
         constructing_unit_Datapath_Middle_registers2_5_n57,
         constructing_unit_Datapath_Middle_registers2_5_n56,
         constructing_unit_Datapath_Middle_registers2_5_n55,
         constructing_unit_Datapath_Middle_registers2_5_n54,
         constructing_unit_Datapath_Middle_registers2_5_n53,
         constructing_unit_Datapath_Middle_registers2_5_n52,
         constructing_unit_Datapath_Middle_registers2_5_n51,
         constructing_unit_Datapath_Middle_registers2_5_n50,
         constructing_unit_Datapath_Middle_registers2_5_n49,
         constructing_unit_Datapath_Middle_registers2_5_n48,
         constructing_unit_Datapath_Middle_registers2_5_n47,
         constructing_unit_Datapath_Middle_registers2_5_n46,
         constructing_unit_Datapath_Middle_registers2_5_n45,
         constructing_unit_Datapath_Middle_registers2_5_n44,
         constructing_unit_Datapath_Middle_registers2_5_n43,
         constructing_unit_Datapath_Middle_registers2_5_n42,
         constructing_unit_Datapath_Middle_registers2_5_n41,
         constructing_unit_Datapath_Middle_registers2_5_n40,
         constructing_unit_Datapath_Middle_registers2_5_n39,
         constructing_unit_Datapath_Middle_registers2_5_n38,
         constructing_unit_Datapath_Middle_registers2_5_n37,
         constructing_unit_Datapath_Middle_registers2_5_n36,
         constructing_unit_Datapath_Middle_registers2_5_n35,
         constructing_unit_Datapath_Middle_registers2_5_n33,
         constructing_unit_Datapath_Middle_registers2_6_n67,
         constructing_unit_Datapath_Middle_registers2_6_n66,
         constructing_unit_Datapath_Middle_registers2_6_n65,
         constructing_unit_Datapath_Middle_registers2_6_n64,
         constructing_unit_Datapath_Middle_registers2_6_n63,
         constructing_unit_Datapath_Middle_registers2_6_n62,
         constructing_unit_Datapath_Middle_registers2_6_n61,
         constructing_unit_Datapath_Middle_registers2_6_n60,
         constructing_unit_Datapath_Middle_registers2_6_n59,
         constructing_unit_Datapath_Middle_registers2_6_n58,
         constructing_unit_Datapath_Middle_registers2_6_n57,
         constructing_unit_Datapath_Middle_registers2_6_n56,
         constructing_unit_Datapath_Middle_registers2_6_n55,
         constructing_unit_Datapath_Middle_registers2_6_n54,
         constructing_unit_Datapath_Middle_registers2_6_n53,
         constructing_unit_Datapath_Middle_registers2_6_n52,
         constructing_unit_Datapath_Middle_registers2_6_n51,
         constructing_unit_Datapath_Middle_registers2_6_n50,
         constructing_unit_Datapath_Middle_registers2_6_n49,
         constructing_unit_Datapath_Middle_registers2_6_n48,
         constructing_unit_Datapath_Middle_registers2_6_n47,
         constructing_unit_Datapath_Middle_registers2_6_n46,
         constructing_unit_Datapath_Middle_registers2_6_n45,
         constructing_unit_Datapath_Middle_registers2_6_n44,
         constructing_unit_Datapath_Middle_registers2_6_n43,
         constructing_unit_Datapath_Middle_registers2_6_n42,
         constructing_unit_Datapath_Middle_registers2_6_n41,
         constructing_unit_Datapath_Middle_registers2_6_n40,
         constructing_unit_Datapath_Middle_registers2_6_n39,
         constructing_unit_Datapath_Middle_registers2_6_n38,
         constructing_unit_Datapath_Middle_registers2_6_n37,
         constructing_unit_Datapath_Middle_registers2_6_n36,
         constructing_unit_Datapath_Middle_registers2_6_n35,
         constructing_unit_Datapath_Middle_registers2_6_n33,
         constructing_unit_Datapath_Middle_registers2_7_n67,
         constructing_unit_Datapath_Middle_registers2_7_n66,
         constructing_unit_Datapath_Middle_registers2_7_n65,
         constructing_unit_Datapath_Middle_registers2_7_n64,
         constructing_unit_Datapath_Middle_registers2_7_n63,
         constructing_unit_Datapath_Middle_registers2_7_n62,
         constructing_unit_Datapath_Middle_registers2_7_n61,
         constructing_unit_Datapath_Middle_registers2_7_n60,
         constructing_unit_Datapath_Middle_registers2_7_n59,
         constructing_unit_Datapath_Middle_registers2_7_n58,
         constructing_unit_Datapath_Middle_registers2_7_n57,
         constructing_unit_Datapath_Middle_registers2_7_n56,
         constructing_unit_Datapath_Middle_registers2_7_n55,
         constructing_unit_Datapath_Middle_registers2_7_n54,
         constructing_unit_Datapath_Middle_registers2_7_n53,
         constructing_unit_Datapath_Middle_registers2_7_n52,
         constructing_unit_Datapath_Middle_registers2_7_n51,
         constructing_unit_Datapath_Middle_registers2_7_n50,
         constructing_unit_Datapath_Middle_registers2_7_n49,
         constructing_unit_Datapath_Middle_registers2_7_n48,
         constructing_unit_Datapath_Middle_registers2_7_n47,
         constructing_unit_Datapath_Middle_registers2_7_n46,
         constructing_unit_Datapath_Middle_registers2_7_n45,
         constructing_unit_Datapath_Middle_registers2_7_n44,
         constructing_unit_Datapath_Middle_registers2_7_n43,
         constructing_unit_Datapath_Middle_registers2_7_n42,
         constructing_unit_Datapath_Middle_registers2_7_n41,
         constructing_unit_Datapath_Middle_registers2_7_n40,
         constructing_unit_Datapath_Middle_registers2_7_n39,
         constructing_unit_Datapath_Middle_registers2_7_n38,
         constructing_unit_Datapath_Middle_registers2_7_n37,
         constructing_unit_Datapath_Middle_registers2_7_n36,
         constructing_unit_Datapath_Middle_registers2_7_n35,
         constructing_unit_Datapath_Middle_registers2_7_n33,
         constructing_unit_Datapath_Middle_registers2_8_n67,
         constructing_unit_Datapath_Middle_registers2_8_n66,
         constructing_unit_Datapath_Middle_registers2_8_n65,
         constructing_unit_Datapath_Middle_registers2_8_n64,
         constructing_unit_Datapath_Middle_registers2_8_n63,
         constructing_unit_Datapath_Middle_registers2_8_n62,
         constructing_unit_Datapath_Middle_registers2_8_n61,
         constructing_unit_Datapath_Middle_registers2_8_n60,
         constructing_unit_Datapath_Middle_registers2_8_n59,
         constructing_unit_Datapath_Middle_registers2_8_n58,
         constructing_unit_Datapath_Middle_registers2_8_n57,
         constructing_unit_Datapath_Middle_registers2_8_n56,
         constructing_unit_Datapath_Middle_registers2_8_n55,
         constructing_unit_Datapath_Middle_registers2_8_n54,
         constructing_unit_Datapath_Middle_registers2_8_n53,
         constructing_unit_Datapath_Middle_registers2_8_n52,
         constructing_unit_Datapath_Middle_registers2_8_n51,
         constructing_unit_Datapath_Middle_registers2_8_n50,
         constructing_unit_Datapath_Middle_registers2_8_n49,
         constructing_unit_Datapath_Middle_registers2_8_n48,
         constructing_unit_Datapath_Middle_registers2_8_n47,
         constructing_unit_Datapath_Middle_registers2_8_n46,
         constructing_unit_Datapath_Middle_registers2_8_n45,
         constructing_unit_Datapath_Middle_registers2_8_n44,
         constructing_unit_Datapath_Middle_registers2_8_n43,
         constructing_unit_Datapath_Middle_registers2_8_n42,
         constructing_unit_Datapath_Middle_registers2_8_n41,
         constructing_unit_Datapath_Middle_registers2_8_n40,
         constructing_unit_Datapath_Middle_registers2_8_n39,
         constructing_unit_Datapath_Middle_registers2_8_n38,
         constructing_unit_Datapath_Middle_registers2_8_n37,
         constructing_unit_Datapath_Middle_registers2_8_n36,
         constructing_unit_Datapath_Middle_registers2_8_n35,
         constructing_unit_Datapath_Middle_registers2_8_n33,
         constructing_unit_Datapath_Middle_registers2_9_n67,
         constructing_unit_Datapath_Middle_registers2_9_n66,
         constructing_unit_Datapath_Middle_registers2_9_n65,
         constructing_unit_Datapath_Middle_registers2_9_n64,
         constructing_unit_Datapath_Middle_registers2_9_n63,
         constructing_unit_Datapath_Middle_registers2_9_n62,
         constructing_unit_Datapath_Middle_registers2_9_n61,
         constructing_unit_Datapath_Middle_registers2_9_n60,
         constructing_unit_Datapath_Middle_registers2_9_n59,
         constructing_unit_Datapath_Middle_registers2_9_n58,
         constructing_unit_Datapath_Middle_registers2_9_n57,
         constructing_unit_Datapath_Middle_registers2_9_n56,
         constructing_unit_Datapath_Middle_registers2_9_n55,
         constructing_unit_Datapath_Middle_registers2_9_n54,
         constructing_unit_Datapath_Middle_registers2_9_n53,
         constructing_unit_Datapath_Middle_registers2_9_n52,
         constructing_unit_Datapath_Middle_registers2_9_n51,
         constructing_unit_Datapath_Middle_registers2_9_n50,
         constructing_unit_Datapath_Middle_registers2_9_n49,
         constructing_unit_Datapath_Middle_registers2_9_n48,
         constructing_unit_Datapath_Middle_registers2_9_n47,
         constructing_unit_Datapath_Middle_registers2_9_n46,
         constructing_unit_Datapath_Middle_registers2_9_n45,
         constructing_unit_Datapath_Middle_registers2_9_n44,
         constructing_unit_Datapath_Middle_registers2_9_n43,
         constructing_unit_Datapath_Middle_registers2_9_n42,
         constructing_unit_Datapath_Middle_registers2_9_n41,
         constructing_unit_Datapath_Middle_registers2_9_n40,
         constructing_unit_Datapath_Middle_registers2_9_n39,
         constructing_unit_Datapath_Middle_registers2_9_n38,
         constructing_unit_Datapath_Middle_registers2_9_n37,
         constructing_unit_Datapath_Middle_registers2_9_n36,
         constructing_unit_Datapath_Middle_registers2_9_n35,
         constructing_unit_Datapath_Middle_registers2_9_n33,
         constructing_unit_Datapath_Middle_registers2_10_n67,
         constructing_unit_Datapath_Middle_registers2_10_n66,
         constructing_unit_Datapath_Middle_registers2_10_n65,
         constructing_unit_Datapath_Middle_registers2_10_n64,
         constructing_unit_Datapath_Middle_registers2_10_n63,
         constructing_unit_Datapath_Middle_registers2_10_n62,
         constructing_unit_Datapath_Middle_registers2_10_n61,
         constructing_unit_Datapath_Middle_registers2_10_n60,
         constructing_unit_Datapath_Middle_registers2_10_n59,
         constructing_unit_Datapath_Middle_registers2_10_n58,
         constructing_unit_Datapath_Middle_registers2_10_n57,
         constructing_unit_Datapath_Middle_registers2_10_n56,
         constructing_unit_Datapath_Middle_registers2_10_n55,
         constructing_unit_Datapath_Middle_registers2_10_n54,
         constructing_unit_Datapath_Middle_registers2_10_n53,
         constructing_unit_Datapath_Middle_registers2_10_n52,
         constructing_unit_Datapath_Middle_registers2_10_n51,
         constructing_unit_Datapath_Middle_registers2_10_n50,
         constructing_unit_Datapath_Middle_registers2_10_n49,
         constructing_unit_Datapath_Middle_registers2_10_n48,
         constructing_unit_Datapath_Middle_registers2_10_n47,
         constructing_unit_Datapath_Middle_registers2_10_n46,
         constructing_unit_Datapath_Middle_registers2_10_n45,
         constructing_unit_Datapath_Middle_registers2_10_n44,
         constructing_unit_Datapath_Middle_registers2_10_n43,
         constructing_unit_Datapath_Middle_registers2_10_n42,
         constructing_unit_Datapath_Middle_registers2_10_n41,
         constructing_unit_Datapath_Middle_registers2_10_n40,
         constructing_unit_Datapath_Middle_registers2_10_n39,
         constructing_unit_Datapath_Middle_registers2_10_n38,
         constructing_unit_Datapath_Middle_registers2_10_n37,
         constructing_unit_Datapath_Middle_registers2_10_n36,
         constructing_unit_Datapath_Middle_registers2_10_n35,
         constructing_unit_Datapath_Middle_registers2_10_n33,
         constructing_unit_Datapath_Middle_registers2_11_n67,
         constructing_unit_Datapath_Middle_registers2_11_n66,
         constructing_unit_Datapath_Middle_registers2_11_n65,
         constructing_unit_Datapath_Middle_registers2_11_n64,
         constructing_unit_Datapath_Middle_registers2_11_n63,
         constructing_unit_Datapath_Middle_registers2_11_n62,
         constructing_unit_Datapath_Middle_registers2_11_n61,
         constructing_unit_Datapath_Middle_registers2_11_n60,
         constructing_unit_Datapath_Middle_registers2_11_n59,
         constructing_unit_Datapath_Middle_registers2_11_n58,
         constructing_unit_Datapath_Middle_registers2_11_n57,
         constructing_unit_Datapath_Middle_registers2_11_n56,
         constructing_unit_Datapath_Middle_registers2_11_n55,
         constructing_unit_Datapath_Middle_registers2_11_n54,
         constructing_unit_Datapath_Middle_registers2_11_n53,
         constructing_unit_Datapath_Middle_registers2_11_n52,
         constructing_unit_Datapath_Middle_registers2_11_n51,
         constructing_unit_Datapath_Middle_registers2_11_n50,
         constructing_unit_Datapath_Middle_registers2_11_n49,
         constructing_unit_Datapath_Middle_registers2_11_n48,
         constructing_unit_Datapath_Middle_registers2_11_n47,
         constructing_unit_Datapath_Middle_registers2_11_n46,
         constructing_unit_Datapath_Middle_registers2_11_n45,
         constructing_unit_Datapath_Middle_registers2_11_n44,
         constructing_unit_Datapath_Middle_registers2_11_n43,
         constructing_unit_Datapath_Middle_registers2_11_n42,
         constructing_unit_Datapath_Middle_registers2_11_n41,
         constructing_unit_Datapath_Middle_registers2_11_n40,
         constructing_unit_Datapath_Middle_registers2_11_n39,
         constructing_unit_Datapath_Middle_registers2_11_n38,
         constructing_unit_Datapath_Middle_registers2_11_n37,
         constructing_unit_Datapath_Middle_registers2_11_n36,
         constructing_unit_Datapath_Middle_registers2_11_n35,
         constructing_unit_Datapath_Middle_registers2_11_n33,
         constructing_unit_Datapath_Middle_registers2_12_n67,
         constructing_unit_Datapath_Middle_registers2_12_n66,
         constructing_unit_Datapath_Middle_registers2_12_n65,
         constructing_unit_Datapath_Middle_registers2_12_n64,
         constructing_unit_Datapath_Middle_registers2_12_n63,
         constructing_unit_Datapath_Middle_registers2_12_n62,
         constructing_unit_Datapath_Middle_registers2_12_n61,
         constructing_unit_Datapath_Middle_registers2_12_n60,
         constructing_unit_Datapath_Middle_registers2_12_n59,
         constructing_unit_Datapath_Middle_registers2_12_n58,
         constructing_unit_Datapath_Middle_registers2_12_n57,
         constructing_unit_Datapath_Middle_registers2_12_n56,
         constructing_unit_Datapath_Middle_registers2_12_n55,
         constructing_unit_Datapath_Middle_registers2_12_n54,
         constructing_unit_Datapath_Middle_registers2_12_n53,
         constructing_unit_Datapath_Middle_registers2_12_n52,
         constructing_unit_Datapath_Middle_registers2_12_n51,
         constructing_unit_Datapath_Middle_registers2_12_n50,
         constructing_unit_Datapath_Middle_registers2_12_n49,
         constructing_unit_Datapath_Middle_registers2_12_n48,
         constructing_unit_Datapath_Middle_registers2_12_n47,
         constructing_unit_Datapath_Middle_registers2_12_n46,
         constructing_unit_Datapath_Middle_registers2_12_n45,
         constructing_unit_Datapath_Middle_registers2_12_n44,
         constructing_unit_Datapath_Middle_registers2_12_n43,
         constructing_unit_Datapath_Middle_registers2_12_n42,
         constructing_unit_Datapath_Middle_registers2_12_n41,
         constructing_unit_Datapath_Middle_registers2_12_n40,
         constructing_unit_Datapath_Middle_registers2_12_n39,
         constructing_unit_Datapath_Middle_registers2_12_n38,
         constructing_unit_Datapath_Middle_registers2_12_n37,
         constructing_unit_Datapath_Middle_registers2_12_n36,
         constructing_unit_Datapath_Middle_registers2_12_n35,
         constructing_unit_Datapath_Middle_registers2_12_n33,
         constructing_unit_Datapath_Middle_registers2_13_n67,
         constructing_unit_Datapath_Middle_registers2_13_n66,
         constructing_unit_Datapath_Middle_registers2_13_n65,
         constructing_unit_Datapath_Middle_registers2_13_n64,
         constructing_unit_Datapath_Middle_registers2_13_n63,
         constructing_unit_Datapath_Middle_registers2_13_n62,
         constructing_unit_Datapath_Middle_registers2_13_n61,
         constructing_unit_Datapath_Middle_registers2_13_n60,
         constructing_unit_Datapath_Middle_registers2_13_n59,
         constructing_unit_Datapath_Middle_registers2_13_n58,
         constructing_unit_Datapath_Middle_registers2_13_n57,
         constructing_unit_Datapath_Middle_registers2_13_n56,
         constructing_unit_Datapath_Middle_registers2_13_n55,
         constructing_unit_Datapath_Middle_registers2_13_n54,
         constructing_unit_Datapath_Middle_registers2_13_n53,
         constructing_unit_Datapath_Middle_registers2_13_n52,
         constructing_unit_Datapath_Middle_registers2_13_n51,
         constructing_unit_Datapath_Middle_registers2_13_n50,
         constructing_unit_Datapath_Middle_registers2_13_n49,
         constructing_unit_Datapath_Middle_registers2_13_n48,
         constructing_unit_Datapath_Middle_registers2_13_n47,
         constructing_unit_Datapath_Middle_registers2_13_n46,
         constructing_unit_Datapath_Middle_registers2_13_n45,
         constructing_unit_Datapath_Middle_registers2_13_n44,
         constructing_unit_Datapath_Middle_registers2_13_n43,
         constructing_unit_Datapath_Middle_registers2_13_n42,
         constructing_unit_Datapath_Middle_registers2_13_n41,
         constructing_unit_Datapath_Middle_registers2_13_n40,
         constructing_unit_Datapath_Middle_registers2_13_n39,
         constructing_unit_Datapath_Middle_registers2_13_n38,
         constructing_unit_Datapath_Middle_registers2_13_n37,
         constructing_unit_Datapath_Middle_registers2_13_n36,
         constructing_unit_Datapath_Middle_registers2_13_n35,
         constructing_unit_Datapath_Middle_registers2_13_n33,
         constructing_unit_Datapath_Last_register0_h_n69,
         constructing_unit_Datapath_Last_register0_h_n68,
         constructing_unit_Datapath_Last_register0_h_n67,
         constructing_unit_Datapath_Last_register0_h_n66,
         constructing_unit_Datapath_Last_register0_h_n65,
         constructing_unit_Datapath_Last_register0_h_n64,
         constructing_unit_Datapath_Last_register0_h_n63,
         constructing_unit_Datapath_Last_register0_h_n62,
         constructing_unit_Datapath_Last_register0_h_n61,
         constructing_unit_Datapath_Last_register0_h_n60,
         constructing_unit_Datapath_Last_register0_h_n59,
         constructing_unit_Datapath_Last_register0_h_n58,
         constructing_unit_Datapath_Last_register0_h_n57,
         constructing_unit_Datapath_Last_register0_h_n56,
         constructing_unit_Datapath_Last_register0_h_n55,
         constructing_unit_Datapath_Last_register0_h_n54,
         constructing_unit_Datapath_Last_register0_h_n53,
         constructing_unit_Datapath_Last_register0_h_n52,
         constructing_unit_Datapath_Last_register0_h_n51,
         constructing_unit_Datapath_Last_register0_h_n50,
         constructing_unit_Datapath_Last_register0_h_n49,
         constructing_unit_Datapath_Last_register0_h_n48,
         constructing_unit_Datapath_Last_register0_h_n47,
         constructing_unit_Datapath_Last_register0_h_n46,
         constructing_unit_Datapath_Last_register0_h_n45,
         constructing_unit_Datapath_Last_register0_h_n44,
         constructing_unit_Datapath_Last_register0_h_n43,
         constructing_unit_Datapath_Last_register0_h_n42,
         constructing_unit_Datapath_Last_register0_h_n41,
         constructing_unit_Datapath_Last_register0_h_n40,
         constructing_unit_Datapath_Last_register0_h_n39,
         constructing_unit_Datapath_Last_register0_h_n38,
         constructing_unit_Datapath_Last_register0_h_n37,
         constructing_unit_Datapath_Last_register0_h_n36,
         constructing_unit_Datapath_Last_register0_h_n35,
         constructing_unit_Datapath_Last_register0_h_n33,
         constructing_unit_Datapath_Last_register1_h_n69,
         constructing_unit_Datapath_Last_register1_h_n68,
         constructing_unit_Datapath_Last_register1_h_n67,
         constructing_unit_Datapath_Last_register1_h_n66,
         constructing_unit_Datapath_Last_register1_h_n65,
         constructing_unit_Datapath_Last_register1_h_n64,
         constructing_unit_Datapath_Last_register1_h_n63,
         constructing_unit_Datapath_Last_register1_h_n62,
         constructing_unit_Datapath_Last_register1_h_n61,
         constructing_unit_Datapath_Last_register1_h_n60,
         constructing_unit_Datapath_Last_register1_h_n59,
         constructing_unit_Datapath_Last_register1_h_n58,
         constructing_unit_Datapath_Last_register1_h_n57,
         constructing_unit_Datapath_Last_register1_h_n56,
         constructing_unit_Datapath_Last_register1_h_n55,
         constructing_unit_Datapath_Last_register1_h_n54,
         constructing_unit_Datapath_Last_register1_h_n53,
         constructing_unit_Datapath_Last_register1_h_n52,
         constructing_unit_Datapath_Last_register1_h_n51,
         constructing_unit_Datapath_Last_register1_h_n50,
         constructing_unit_Datapath_Last_register1_h_n49,
         constructing_unit_Datapath_Last_register1_h_n48,
         constructing_unit_Datapath_Last_register1_h_n47,
         constructing_unit_Datapath_Last_register1_h_n46,
         constructing_unit_Datapath_Last_register1_h_n45,
         constructing_unit_Datapath_Last_register1_h_n44,
         constructing_unit_Datapath_Last_register1_h_n43,
         constructing_unit_Datapath_Last_register1_h_n42,
         constructing_unit_Datapath_Last_register1_h_n41,
         constructing_unit_Datapath_Last_register1_h_n40,
         constructing_unit_Datapath_Last_register1_h_n39,
         constructing_unit_Datapath_Last_register1_h_n38,
         constructing_unit_Datapath_Last_register1_h_n37,
         constructing_unit_Datapath_Last_register1_h_n36,
         constructing_unit_Datapath_Last_register1_h_n35,
         constructing_unit_Datapath_Last_register1_h_n33,
         constructing_unit_Datapath_Last_register2_h_n69,
         constructing_unit_Datapath_Last_register2_h_n68,
         constructing_unit_Datapath_Last_register2_h_n67,
         constructing_unit_Datapath_Last_register2_h_n66,
         constructing_unit_Datapath_Last_register2_h_n65,
         constructing_unit_Datapath_Last_register2_h_n64,
         constructing_unit_Datapath_Last_register2_h_n63,
         constructing_unit_Datapath_Last_register2_h_n62,
         constructing_unit_Datapath_Last_register2_h_n61,
         constructing_unit_Datapath_Last_register2_h_n60,
         constructing_unit_Datapath_Last_register2_h_n59,
         constructing_unit_Datapath_Last_register2_h_n58,
         constructing_unit_Datapath_Last_register2_h_n57,
         constructing_unit_Datapath_Last_register2_h_n56,
         constructing_unit_Datapath_Last_register2_h_n55,
         constructing_unit_Datapath_Last_register2_h_n54,
         constructing_unit_Datapath_Last_register2_h_n53,
         constructing_unit_Datapath_Last_register2_h_n52,
         constructing_unit_Datapath_Last_register2_h_n51,
         constructing_unit_Datapath_Last_register2_h_n50,
         constructing_unit_Datapath_Last_register2_h_n49,
         constructing_unit_Datapath_Last_register2_h_n48,
         constructing_unit_Datapath_Last_register2_h_n47,
         constructing_unit_Datapath_Last_register2_h_n46,
         constructing_unit_Datapath_Last_register2_h_n45,
         constructing_unit_Datapath_Last_register2_h_n44,
         constructing_unit_Datapath_Last_register2_h_n43,
         constructing_unit_Datapath_Last_register2_h_n42,
         constructing_unit_Datapath_Last_register2_h_n41,
         constructing_unit_Datapath_Last_register2_h_n40,
         constructing_unit_Datapath_Last_register2_h_n39,
         constructing_unit_Datapath_Last_register2_h_n38,
         constructing_unit_Datapath_Last_register2_h_n37,
         constructing_unit_Datapath_Last_register2_h_n36,
         constructing_unit_Datapath_Last_register2_h_n35,
         constructing_unit_Datapath_Last_register2_h_n33,
         extimating_unit_SAD_tmp_RST_CU_int, extimating_unit_LE_ab_CU_int,
         extimating_unit_READY_RST_int, extimating_unit_RST2_int,
         extimating_unit_RST1_int, extimating_unit_RST_BLKy_int,
         extimating_unit_CE_BLKy_int, extimating_unit_CE_REPy_int,
         extimating_unit_RST_BLKx_int, extimating_unit_CE_BLKx_int,
         extimating_unit_CE_REPx_int, extimating_unit_RF_in_WE_int,
         extimating_unit_RF_Addr_DP_int, extimating_unit_VALID_int,
         extimating_unit_Pixel_Retrieval_Unit_n130,
         extimating_unit_Pixel_Retrieval_Unit_n129,
         extimating_unit_Pixel_Retrieval_Unit_n128,
         extimating_unit_Pixel_Retrieval_Unit_n127,
         extimating_unit_Pixel_Retrieval_Unit_n126,
         extimating_unit_Pixel_Retrieval_Unit_n125,
         extimating_unit_Pixel_Retrieval_Unit_n124,
         extimating_unit_Pixel_Retrieval_Unit_n123,
         extimating_unit_Pixel_Retrieval_Unit_n122,
         extimating_unit_Pixel_Retrieval_Unit_n121,
         extimating_unit_Pixel_Retrieval_Unit_n120,
         extimating_unit_Pixel_Retrieval_Unit_n119,
         extimating_unit_Pixel_Retrieval_Unit_n118,
         extimating_unit_Pixel_Retrieval_Unit_n117,
         extimating_unit_Pixel_Retrieval_Unit_n116,
         extimating_unit_Pixel_Retrieval_Unit_n115,
         extimating_unit_Pixel_Retrieval_Unit_n114,
         extimating_unit_Pixel_Retrieval_Unit_n113,
         extimating_unit_Pixel_Retrieval_Unit_n112,
         extimating_unit_Pixel_Retrieval_Unit_n111,
         extimating_unit_Pixel_Retrieval_Unit_n110,
         extimating_unit_Pixel_Retrieval_Unit_n109,
         extimating_unit_Pixel_Retrieval_Unit_n108,
         extimating_unit_Pixel_Retrieval_Unit_n107,
         extimating_unit_Pixel_Retrieval_Unit_n106,
         extimating_unit_Pixel_Retrieval_Unit_n105,
         extimating_unit_Pixel_Retrieval_Unit_n104,
         extimating_unit_Pixel_Retrieval_Unit_n103,
         extimating_unit_Pixel_Retrieval_Unit_n102,
         extimating_unit_Pixel_Retrieval_Unit_n101,
         extimating_unit_Pixel_Retrieval_Unit_n100,
         extimating_unit_Pixel_Retrieval_Unit_n99,
         extimating_unit_Pixel_Retrieval_Unit_n74,
         extimating_unit_Pixel_Retrieval_Unit_n73,
         extimating_unit_Pixel_Retrieval_Unit_n72,
         extimating_unit_Pixel_Retrieval_Unit_n71,
         extimating_unit_Pixel_Retrieval_Unit_n70,
         extimating_unit_Pixel_Retrieval_Unit_n69,
         extimating_unit_Pixel_Retrieval_Unit_n68,
         extimating_unit_Pixel_Retrieval_Unit_n67,
         extimating_unit_Pixel_Retrieval_Unit_n66,
         extimating_unit_Pixel_Retrieval_Unit_n65,
         extimating_unit_Pixel_Retrieval_Unit_n64,
         extimating_unit_Pixel_Retrieval_Unit_n63,
         extimating_unit_Pixel_Retrieval_Unit_n62,
         extimating_unit_Pixel_Retrieval_Unit_n61,
         extimating_unit_Pixel_Retrieval_Unit_n60,
         extimating_unit_Pixel_Retrieval_Unit_n59,
         extimating_unit_Pixel_Retrieval_Unit_n58,
         extimating_unit_Pixel_Retrieval_Unit_n57,
         extimating_unit_Pixel_Retrieval_Unit_n56,
         extimating_unit_Pixel_Retrieval_Unit_n55,
         extimating_unit_Pixel_Retrieval_Unit_n54,
         extimating_unit_Pixel_Retrieval_Unit_n53,
         extimating_unit_Pixel_Retrieval_Unit_n52,
         extimating_unit_Pixel_Retrieval_Unit_n51,
         extimating_unit_Pixel_Retrieval_Unit_n50,
         extimating_unit_Pixel_Retrieval_Unit_n49,
         extimating_unit_Pixel_Retrieval_Unit_n48,
         extimating_unit_Pixel_Retrieval_Unit_n47,
         extimating_unit_Pixel_Retrieval_Unit_n46,
         extimating_unit_Pixel_Retrieval_Unit_n45,
         extimating_unit_Pixel_Retrieval_Unit_n44,
         extimating_unit_Pixel_Retrieval_Unit_n43,
         extimating_unit_Pixel_Retrieval_Unit_n42,
         extimating_unit_Pixel_Retrieval_Unit_n41,
         extimating_unit_Pixel_Retrieval_Unit_n40,
         extimating_unit_Pixel_Retrieval_Unit_n39,
         extimating_unit_Pixel_Retrieval_Unit_n38,
         extimating_unit_Pixel_Retrieval_Unit_n37,
         extimating_unit_Pixel_Retrieval_Unit_n36,
         extimating_unit_Pixel_Retrieval_Unit_n35,
         extimating_unit_Pixel_Retrieval_Unit_n34,
         extimating_unit_Pixel_Retrieval_Unit_n33,
         extimating_unit_Pixel_Retrieval_Unit_n32,
         extimating_unit_Pixel_Retrieval_Unit_n31,
         extimating_unit_Pixel_Retrieval_Unit_n30,
         extimating_unit_Pixel_Retrieval_Unit_n29,
         extimating_unit_Pixel_Retrieval_Unit_n28,
         extimating_unit_Pixel_Retrieval_Unit_n27,
         extimating_unit_Pixel_Retrieval_Unit_n26,
         extimating_unit_Pixel_Retrieval_Unit_n25,
         extimating_unit_Pixel_Retrieval_Unit_n24,
         extimating_unit_Pixel_Retrieval_Unit_n23,
         extimating_unit_Pixel_Retrieval_Unit_n22,
         extimating_unit_Pixel_Retrieval_Unit_n21,
         extimating_unit_Pixel_Retrieval_Unit_n20,
         extimating_unit_Pixel_Retrieval_Unit_n19,
         extimating_unit_Pixel_Retrieval_Unit_n18,
         extimating_unit_Pixel_Retrieval_Unit_n17,
         extimating_unit_Pixel_Retrieval_Unit_n16,
         extimating_unit_Pixel_Retrieval_Unit_n15,
         extimating_unit_Pixel_Retrieval_Unit_n14,
         extimating_unit_Pixel_Retrieval_Unit_n13,
         extimating_unit_Pixel_Retrieval_Unit_n12,
         extimating_unit_Pixel_Retrieval_Unit_n11,
         extimating_unit_Pixel_Retrieval_Unit_n9,
         extimating_unit_Pixel_Retrieval_Unit_n8,
         extimating_unit_Pixel_Retrieval_Unit_n7,
         extimating_unit_Pixel_Retrieval_Unit_n6,
         extimating_unit_Pixel_Retrieval_Unit_n5,
         extimating_unit_Pixel_Retrieval_Unit_n4,
         extimating_unit_Pixel_Retrieval_Unit_n3,
         extimating_unit_Pixel_Retrieval_Unit_n2,
         extimating_unit_Pixel_Retrieval_Unit_n1,
         extimating_unit_Pixel_Retrieval_Unit_add_239_carry_2_,
         extimating_unit_Pixel_Retrieval_Unit_n98,
         extimating_unit_Pixel_Retrieval_Unit_n97,
         extimating_unit_Pixel_Retrieval_Unit_n96,
         extimating_unit_Pixel_Retrieval_Unit_n95,
         extimating_unit_Pixel_Retrieval_Unit_n94,
         extimating_unit_Pixel_Retrieval_Unit_n93,
         extimating_unit_Pixel_Retrieval_Unit_n92,
         extimating_unit_Pixel_Retrieval_Unit_n91,
         extimating_unit_Pixel_Retrieval_Unit_n90,
         extimating_unit_Pixel_Retrieval_Unit_n89,
         extimating_unit_Pixel_Retrieval_Unit_n88,
         extimating_unit_Pixel_Retrieval_Unit_n87,
         extimating_unit_Pixel_Retrieval_Unit_n86,
         extimating_unit_Pixel_Retrieval_Unit_n85,
         extimating_unit_Pixel_Retrieval_Unit_n84,
         extimating_unit_Pixel_Retrieval_Unit_n83,
         extimating_unit_Pixel_Retrieval_Unit_n82,
         extimating_unit_Pixel_Retrieval_Unit_n81,
         extimating_unit_Pixel_Retrieval_Unit_n80,
         extimating_unit_Pixel_Retrieval_Unit_n79,
         extimating_unit_Pixel_Retrieval_Unit_n78,
         extimating_unit_Pixel_Retrieval_Unit_n77,
         extimating_unit_Pixel_Retrieval_Unit_n76,
         extimating_unit_Pixel_Retrieval_Unit_n75,
         extimating_unit_Pixel_Retrieval_Unit_y_short_1_,
         extimating_unit_Pixel_Retrieval_Unit_y_count_out_0_,
         extimating_unit_Pixel_Retrieval_Unit_y_count_out_1_,
         extimating_unit_Pixel_Retrieval_Unit_x_0_,
         extimating_unit_Pixel_Retrieval_Unit_x_1_,
         extimating_unit_Pixel_Retrieval_Unit_x_2_,
         extimating_unit_Pixel_Retrieval_Unit_x_3_,
         extimating_unit_Pixel_Retrieval_Unit_x_4_,
         extimating_unit_Pixel_Retrieval_Unit_x_5_,
         extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__0_,
         extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__1_,
         extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__2_,
         extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__3_,
         extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__4_,
         extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__5_,
         extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__0_,
         extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__1_,
         extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__2_,
         extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__3_,
         extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__4_,
         extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__5_,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__0_,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__1_,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__2_,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__3_,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__4_,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__5_,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__6_,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__7_,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__8_,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__9_,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__10_,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__11_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__0_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__1_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__2_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__3_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__4_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__5_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__6_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__7_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__8_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__9_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__10_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__0_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__1_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__2_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__3_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__4_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__5_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__6_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__7_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__8_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__9_,
         extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__10_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_0__3_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_0__4_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_0__5_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_1__0_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_1__1_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_1__2_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_1__3_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_1__4_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_1__5_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_2__0_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_2__1_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_2__2_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_2__3_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_2__4_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_2__5_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_3__0_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_3__1_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_3__2_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_3__3_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_3__4_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_3__5_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_5__0_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_5__1_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_5__2_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_5__3_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_5__4_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_5__5_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_6__0_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_6__1_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_6__2_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_6__3_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_6__4_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_6__5_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_7__0_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_7__1_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_7__2_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_7__3_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_7__4_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_7__5_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_8__0_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_8__1_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_8__2_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_8__3_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_8__4_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_8__5_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_9__0_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_9__1_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_9__2_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_9__3_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_9__4_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_9__5_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_10__0_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_10__1_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_10__2_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_10__3_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_10__4_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_10__5_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_11__0_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_11__1_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_11__2_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_11__3_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_11__4_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_11__5_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_12__0_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_12__1_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_12__2_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_12__3_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_12__4_,
         extimating_unit_Pixel_Retrieval_Unit_y0_int_12__5_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_0__3_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_0__4_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_0__5_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_1__0_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_1__1_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_1__2_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_1__3_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_1__4_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_1__5_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_2__0_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_2__1_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_2__2_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_2__3_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_2__4_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_2__5_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_3__0_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_3__1_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_3__2_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_3__3_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_3__4_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_3__5_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_5__0_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_5__1_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_5__2_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_5__3_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_5__4_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_5__5_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_6__0_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_6__1_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_6__2_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_6__3_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_6__4_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_6__5_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_7__0_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_7__1_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_7__2_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_7__3_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_7__4_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_7__5_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_8__0_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_8__1_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_8__2_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_8__3_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_8__4_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_8__5_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_9__0_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_9__1_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_9__2_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_9__3_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_9__4_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_9__5_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_10__0_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_10__1_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_10__2_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_10__3_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_10__4_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_10__5_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_11__0_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_11__1_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_11__2_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_11__3_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_11__4_,
         extimating_unit_Pixel_Retrieval_Unit_x0_int_11__5_,
         extimating_unit_Pixel_Retrieval_Unit_sixPar_samp,
         extimating_unit_Pixel_Retrieval_Unit_CurCU_h_short_0_,
         extimating_unit_Pixel_Retrieval_Unit_CurCU_w_short_0_,
         extimating_unit_Pixel_Retrieval_Unit_width_register_n1,
         extimating_unit_Pixel_Retrieval_Unit_height_register_n1,
         extimating_unit_Pixel_Retrieval_Unit_sixPar_reg_n1,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n416,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n415,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n414,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n413,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n412,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n411,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n410,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n409,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n408,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n407,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n406,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n405,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n404,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n403,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n402,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n401,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n400,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n399,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n398,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n397,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n396,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n395,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n394,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n393,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n392,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n391,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n390,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n389,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n388,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n387,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n386,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n385,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n384,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n383,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n382,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n381,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n380,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n379,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n378,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n377,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n376,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n375,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n374,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n373,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n372,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n371,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n370,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n369,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n368,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n367,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n366,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n365,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n364,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n363,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n362,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n361,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n360,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n359,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n358,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n357,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n356,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n355,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n354,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n353,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n352,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n351,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n350,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n349,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n348,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n347,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n346,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n345,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n344,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n343,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n342,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n341,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n340,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n339,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n338,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n336,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n72,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n71,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n70,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n69,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n68,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n67,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n66,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n65,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n64,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n63,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n62,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n61,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n60,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n59,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n58,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n57,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n56,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n55,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n54,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n53,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n52,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n51,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n50,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n49,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n48,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n47,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n46,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n45,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n44,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n43,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n42,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n41,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n40,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n39,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n38,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n37,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n36,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n35,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n34,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n33,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n32,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n31,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n30,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n29,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n28,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n27,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n26,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n25,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n24,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n23,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n22,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n21,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n20,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n19,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n18,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n17,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n16,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n15,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n13,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n12,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n11,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n10,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n9,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n8,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n7,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n6,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n5,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n4,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n3,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n2,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n337,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n335,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n334,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n333,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n332,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n331,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n330,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n329,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n328,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n327,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n326,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n325,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n324,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n323,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n322,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n321,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n320,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n319,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n318,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n317,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n316,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n315,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n314,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n313,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n312,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n311,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n310,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n309,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n308,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n307,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n306,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n305,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n304,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n303,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n302,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n301,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n300,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n299,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n298,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n297,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n296,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n295,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n294,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n293,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n292,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n291,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n290,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n289,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n288,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n287,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n286,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n285,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n284,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n283,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n282,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n281,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n280,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n279,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n278,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n277,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n276,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n275,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n274,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n273,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n272,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n271,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n270,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n269,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n268,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n267,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n266,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n265,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n264,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n263,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n262,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n261,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n260,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n259,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n258,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n257,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n256,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n255,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n254,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n253,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n252,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n251,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n250,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n249,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n248,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n247,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n246,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n245,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n244,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n243,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n242,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n241,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n240,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n239,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n238,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n237,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n236,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n235,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n234,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n233,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n232,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n231,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n230,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n229,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n228,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n227,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n226,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n225,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n224,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n223,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n222,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n221,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n220,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n219,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n218,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n217,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n216,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n215,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n214,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n213,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n212,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n211,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n210,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n209,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n208,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n207,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n206,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n205,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n204,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n203,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n202,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n201,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n200,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n199,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n198,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n197,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n196,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n195,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n194,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n193,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n192,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n191,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n190,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n189,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n188,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n187,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n186,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n185,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n184,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n183,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n182,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n181,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n180,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n179,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n178,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n177,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n176,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n175,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n174,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n173,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n172,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n171,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n170,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n169,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n168,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n167,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n166,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n165,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n164,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n163,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n162,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n161,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n160,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n159,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n158,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n157,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n156,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n155,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n154,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n153,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n152,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n151,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n150,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n149,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n148,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n147,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n146,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n145,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n144,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n143,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n142,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n141,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n140,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n139,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n138,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n137,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n136,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n135,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n134,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n133,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n132,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n131,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n130,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n129,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n128,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n127,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n126,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n125,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n124,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n123,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n122,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n121,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n120,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n119,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n118,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n117,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n116,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n115,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n114,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n113,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n112,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n111,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n110,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n109,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n108,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n107,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n106,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n105,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n104,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n103,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n102,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n101,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n100,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n99,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n98,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n97,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n96,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n95,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n94,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n93,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n92,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n91,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n90,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n89,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n88,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n87,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n86,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n85,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n84,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n83,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n82,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n81,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n80,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n79,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n78,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n77,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n76,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n75,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n74,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n73,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n14,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_n1,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_samp,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_n7,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_n6,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_n5,
         extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_n3,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_n2,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_n1,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_count_RST,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurRep_n1,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurRep_n2,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n5,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n4,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n3,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n2,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n1,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_n4,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_n3,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_count_RST,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurRep_n3,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurRep_n1,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n10,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n9,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n8,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n7,
         extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n6,
         extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_n1,
         extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_n1,
         extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_n1,
         extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_n1,
         extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_n1,
         extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_n1,
         extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_n1,
         extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_n1,
         extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_n1,
         extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_n1,
         extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_n1,
         extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_n1,
         extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_n1,
         extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_n1,
         extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_n1,
         extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_n1,
         extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_n1,
         extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_n1,
         extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_n1,
         extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_n1,
         extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_n1,
         extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_n1,
         extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_n1,
         extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_n1,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n12,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n11,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n10,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n9,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n8,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n7,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n6,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n5,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n4,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n3,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n2,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n1,
         extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_0_n1,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n12,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n11,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n10,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n9,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n8,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n7,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n6,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n5,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n4,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n3,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n2,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n1,
         extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_1_n1,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n12,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n11,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n10,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n9,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n8,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n7,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n6,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n5,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n4,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n3,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n2,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n1,
         extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_2_n1,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n12,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n11,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n10,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n9,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n8,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n7,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n6,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n5,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n4,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n3,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n2,
         extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n1,
         extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_3_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_en2,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_en1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n65,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n64,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n62,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n61,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n60,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n59,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n58,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n57,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n56,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n55,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n54,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n53,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n52,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n51,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n50,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n49,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n48,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n47,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n46,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n45,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n44,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n43,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n42,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n41,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n16,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n15,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n14,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n13,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n12,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n11,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n10,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n9,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n8,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n7,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n6,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n5,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n4,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n2,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_en2_gen_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n65,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n64,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n62,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n61,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n60,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n59,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n58,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n57,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n56,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n55,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n54,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n53,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n52,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n51,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n50,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n49,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n48,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n47,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n46,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n45,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n44,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n43,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n42,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n41,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n16,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n15,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n14,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n13,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n12,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n11,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n10,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n9,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n8,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n7,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n6,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n5,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n4,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n2,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_en2,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_en1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n65,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n64,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n62,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n61,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n60,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n59,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n58,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n57,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n56,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n55,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n54,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n53,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n52,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n51,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n50,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n49,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n48,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n47,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n46,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n45,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n44,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n43,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n42,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n41,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n16,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n15,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n14,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n13,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n12,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n11,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n10,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n9,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n8,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n7,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n6,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n5,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n4,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n2,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_en2_gen_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n65,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n64,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n62,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n61,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n60,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n59,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n58,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n57,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n56,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n55,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n54,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n53,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n52,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n51,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n50,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n49,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n48,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n47,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n46,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n45,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n44,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n43,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n42,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n41,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n16,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n15,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n14,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n13,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n12,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n11,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n10,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n9,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n8,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n7,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n6,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n5,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n4,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n2,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_en2,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_en1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n65,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n64,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n62,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n61,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n60,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n59,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n58,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n57,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n56,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n55,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n54,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n53,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n52,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n51,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n50,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n49,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n48,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n47,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n46,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n45,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n44,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n43,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n42,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n41,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n16,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n15,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n14,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n13,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n12,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n11,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n10,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n9,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n8,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n7,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n6,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n5,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n4,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n2,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_en2_gen_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n65,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n64,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n62,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n61,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n60,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n59,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n58,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n57,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n56,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n55,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n54,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n53,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n52,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n51,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n50,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n49,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n48,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n47,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n46,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n45,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n44,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n43,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n42,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n41,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n16,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n15,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n14,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n13,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n12,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n11,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n10,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n9,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n8,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n7,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n6,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n5,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n4,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n2,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_en2,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_en1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n65,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n64,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n62,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n61,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n60,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n59,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n58,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n57,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n56,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n55,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n54,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n53,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n52,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n51,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n50,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n49,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n48,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n47,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n46,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n45,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n44,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n43,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n42,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n41,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n16,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n15,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n14,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n13,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n12,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n11,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n10,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n9,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n8,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n7,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n6,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n5,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n4,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n2,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_en2_gen_n1,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n65,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n64,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n62,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n61,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n60,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n59,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n58,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n57,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n56,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n55,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n54,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n53,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n52,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n51,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n50,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n49,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n48,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n47,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n46,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n45,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n44,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n43,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n42,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n41,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n16,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n15,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n14,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n13,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n12,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n11,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n10,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n9,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n8,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n7,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n6,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n5,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n4,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n2,
         extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n37,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n35,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n34,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n33,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n32,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n31,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n30,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n29,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n28,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n27,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n26,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n25,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n24,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n23,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n22,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n21,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n20,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n19,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n18,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n17,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n16,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n15,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n14,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n13,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n12,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n11,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n10,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n9,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n8,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n7,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n6,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n5,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n4,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n3,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n2,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n1,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n75,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n74,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n73,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n72,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n71,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n70,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n69,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n68,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n67,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n66,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n65,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n64,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n63,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n62,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n61,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n60,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n59,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n58,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n57,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n56,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n55,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n54,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n53,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n52,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n51,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n50,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n49,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n48,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n47,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n46,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n45,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n44,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n43,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n42,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n41,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n40,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n75,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n74,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n73,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n72,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n71,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n70,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n69,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n68,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n67,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n66,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n65,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n64,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n63,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n62,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n61,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n60,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n59,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n58,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n57,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n56,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n55,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n54,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n53,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n52,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n51,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n50,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n49,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n48,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n47,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n46,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n45,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n44,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n43,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n42,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n41,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n40,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n75,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n74,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n73,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n72,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n71,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n70,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n69,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n68,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n67,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n66,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n65,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n64,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n63,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n62,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n61,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n60,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n59,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n58,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n57,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n56,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n55,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n54,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n53,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n52,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n51,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n50,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n49,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n48,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n47,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n46,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n45,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n44,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n43,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n42,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n41,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n40,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38,
         extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n41,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n40,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n39,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n38,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n37,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n36,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n35,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n34,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n32,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n31,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n30,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n29,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n28,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n27,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n26,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n25,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n24,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n23,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n22,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n21,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n20,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n19,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n18,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n17,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n16,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n15,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n14,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n13,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n12,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n11,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n10,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n9,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n8,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n7,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n6,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n5,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n4,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n3,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n99,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n98,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n97,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n96,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n95,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n94,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n93,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n92,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n91,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n90,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n89,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n88,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n87,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n86,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n85,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n84,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n83,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n82,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n81,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n80,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n79,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n78,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n77,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n76,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n75,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n73,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n72,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n71,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n70,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n69,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n68,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n67,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n66,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n65,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n64,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n63,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n62,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n61,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n60,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n59,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n58,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n56,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n54,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n53,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n52,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n51,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n50,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n49,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n48,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n47,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n46,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n45,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n44,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n43,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n42,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_result_LE,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_N35,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_2_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_3_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_4_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_5_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_7_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_8_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_9_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_10_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_11_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_12_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_13_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_14_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_15_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_16_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_17_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_18_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_19_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_20_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_21_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_22_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_23_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_24_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_25_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_rst_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_rst_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_int_LE,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_2_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_3_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_4_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_5_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_7_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_8_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_9_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_10_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_11_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_12_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op2_int_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op1_int_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_18_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_19_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_20_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_21_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_22_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_23_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n7,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n5,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n4,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n3,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_SUM_14_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_int_LE_FF_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_RST_FFX_1_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_RST_FFX_2_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_RST_FFX_2_Q,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_result_LE_FF_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n74,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n72,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n73,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n71,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n70,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n69,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n68,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n67,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n66,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n65,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n64,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n63,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n62,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n61,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n60,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n59,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n58,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n57,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n56,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n55,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n54,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n53,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n52,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n51,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n50,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n49,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n48,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n47,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n46,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n45,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n44,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n43,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n42,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n41,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n40,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n39,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n38,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n37,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n36,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n35,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n34,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n33,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n32,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n31,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n30,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n29,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n28,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n27,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n26,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n25,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n24,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n23,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n22,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n21,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n20,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n19,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n18,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n17,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n16,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n15,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n14,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n13,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n12,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n11,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n10,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n9,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n8,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n7,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n6,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n5,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n4,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n3,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n181,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n180,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n179,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n178,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n177,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n176,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n175,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n174,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n173,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n172,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n171,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n170,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n169,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n168,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n120,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n119,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n118,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n117,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n116,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n115,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n114,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n113,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n112,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n111,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n110,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n109,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n108,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n107,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n106,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n105,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n104,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n103,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n102,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n101,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n100,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n99,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n98,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n97,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n95,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n94,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n93,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n92,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n91,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n90,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n89,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n88,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n87,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n86,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n85,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n83,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n82,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n81,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n80,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n79,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n78,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n77,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n76,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n75,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n74,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n73,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n72,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n71,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n70,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n69,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n68,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n67,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n66,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n65,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n64,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n63,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n62,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n61,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n60,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n59,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n58,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n57,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n56,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n55,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n54,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n53,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n52,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n51,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n50,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n49,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n48,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n47,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n46,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n45,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n44,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n43,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n42,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n41,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n40,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n39,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n38,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n37,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n36,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n35,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n34,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n33,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n32,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n31,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n30,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n29,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n28,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n27,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n26,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n25,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n24,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n23,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n22,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n21,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n20,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n19,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n18,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n17,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n16,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n15,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n14,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n13,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n12,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n11,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n10,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n9,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n8,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n7,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n6,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n5,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n4,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n3,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n157,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n156,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n155,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n154,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n153,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n152,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n151,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n150,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n149,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n148,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n147,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n146,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n145,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n143,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n141,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n140,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n139,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n138,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n137,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n136,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n135,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n134,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n133,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n132,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n131,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n130,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n129,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n128,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n127,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n126,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n124,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n123,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n122,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n121,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n120,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n119,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n118,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n117,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n116,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n115,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n114,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n113,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n112,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n111,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n110,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n109,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n108,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n107,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n106,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n105,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n104,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n103,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n102,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n101,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n100,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n41,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n40,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n39,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n38,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n37,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n36,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n35,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n33,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n32,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n31,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n30,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n29,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n28,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n27,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n26,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n25,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n24,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n23,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n22,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n21,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n20,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n19,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n18,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n17,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n16,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n15,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n14,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n13,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n12,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n11,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n10,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n9,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n8,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n7,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n6,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n5,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n4,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n3,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_result_LE,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_N35,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_2_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_3_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_4_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_5_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_7_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_8_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_9_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_10_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_11_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_12_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_13_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_14_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_15_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_16_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_17_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_18_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_19_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_20_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_21_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_22_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_23_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_24_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_25_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_rst_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_rst_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_int_LE,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_2_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_3_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_4_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_5_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_7_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_8_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_9_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_10_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_11_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_12_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op2_int_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op1_int_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_18_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_19_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_20_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_21_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_22_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_23_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n10,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n9,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n8,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n7,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n6,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_SUM_14_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_int_LE_FF_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_RST_FFX_1_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_RST_FFX_2_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_RST_FFX_2_Q,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_result_LE_FF_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n152,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n151,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n150,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n149,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n148,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n147,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n146,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n145,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n144,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n143,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n142,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n141,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n140,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n139,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n138,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n137,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n136,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n135,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n134,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n133,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n132,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n131,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n130,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n129,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n128,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n127,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n126,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n125,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n124,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n123,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n122,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n121,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n120,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n119,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n118,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n117,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n116,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n115,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n114,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n113,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n112,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n111,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n110,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n109,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n108,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n107,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n106,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n105,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n104,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n103,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n102,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n101,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n100,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n99,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n98,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n97,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n96,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n95,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n94,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n93,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n92,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n91,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n90,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n89,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n88,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n87,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n86,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n85,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n84,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n83,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n82,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n81,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n74,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n72,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n181,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n180,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n179,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n178,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n177,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n176,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n175,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n174,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n173,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n172,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n171,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n170,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n169,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n168,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n120,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n119,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n118,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n117,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n116,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n115,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n114,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n113,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n112,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n111,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n110,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n109,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n108,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n107,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n106,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n105,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n104,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n103,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n102,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n101,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n100,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n99,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n98,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n97,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n95,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n94,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n93,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n92,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n91,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n90,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n89,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n88,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n87,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n86,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n85,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n83,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n82,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n81,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n80,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n79,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n78,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n77,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n76,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n75,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n74,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n73,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n72,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n71,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n70,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n69,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n68,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n67,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n66,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n65,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n64,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n63,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n62,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n61,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n60,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n59,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n58,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n57,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n56,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n55,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n54,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n53,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n52,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n51,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n50,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n49,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n48,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n47,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n46,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n45,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n44,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n43,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n42,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n41,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n40,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n39,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n38,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n37,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n36,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n35,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n34,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n33,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n32,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n31,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n30,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n29,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n28,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n27,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n26,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n25,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n24,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n23,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n22,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n21,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n20,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n19,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n18,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n17,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n16,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n15,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n14,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n13,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n12,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n11,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n10,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n9,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n8,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n7,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n6,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n5,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n4,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n3,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n157,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n156,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n155,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n154,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n153,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n152,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n151,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n150,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n149,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n148,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n147,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n146,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n145,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n143,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n141,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n140,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n139,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n138,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n137,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n136,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n135,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n134,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n133,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n132,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n131,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n130,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n129,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n128,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n127,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n126,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n124,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n123,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n122,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n121,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n120,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n119,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n118,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n117,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n116,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n115,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n114,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n113,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n112,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n111,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n110,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n109,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n108,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n107,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n106,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n105,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n104,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n103,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n102,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n101,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n100,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n41,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n40,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n39,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n38,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n37,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n36,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n35,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n33,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n32,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n31,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n30,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n29,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n28,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n27,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n26,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n25,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n24,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n23,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n22,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n21,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n20,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n19,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n18,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n17,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n16,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n15,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n14,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n13,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n12,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n11,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n10,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n9,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n8,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n7,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n6,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n5,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n4,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n3,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_result_LE,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_N35,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_2_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_3_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_4_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_5_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_7_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_8_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_9_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_10_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_11_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_12_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_13_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_14_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_15_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_16_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_17_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_18_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_19_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_20_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_21_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_22_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_23_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_24_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_25_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_rst_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_rst_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_int_LE,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_2_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_3_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_4_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_5_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_7_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_8_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_9_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_10_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_11_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_12_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op2_int_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op1_int_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_18_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_19_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_20_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_21_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_22_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_23_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n10,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n9,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n8,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n7,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n6,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_SUM_14_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_int_LE_FF_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_RST_FFX_1_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_RST_FFX_2_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_RST_FFX_2_Q,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_result_LE_FF_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n152,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n151,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n150,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n149,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n148,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n147,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n146,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n145,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n144,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n143,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n142,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n141,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n140,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n139,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n138,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n137,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n136,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n135,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n134,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n133,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n132,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n131,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n130,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n129,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n128,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n127,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n126,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n125,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n124,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n123,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n122,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n121,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n120,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n119,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n118,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n117,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n116,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n115,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n114,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n113,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n112,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n111,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n110,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n109,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n108,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n107,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n106,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n105,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n104,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n103,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n102,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n101,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n100,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n99,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n98,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n97,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n96,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n95,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n94,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n93,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n92,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n91,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n90,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n89,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n88,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n87,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n86,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n85,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n84,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n83,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n82,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n81,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n74,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n72,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n181,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n180,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n179,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n178,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n177,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n176,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n175,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n174,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n173,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n172,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n171,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n170,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n169,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n168,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n120,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n119,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n118,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n117,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n116,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n115,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n114,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n113,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n112,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n111,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n110,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n109,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n108,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n107,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n106,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n105,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n104,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n103,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n102,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n101,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n100,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n99,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n98,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n97,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n95,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n94,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n93,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n92,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n91,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n90,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n89,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n88,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n87,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n86,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n85,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n83,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n82,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n81,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n80,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n79,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n78,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n77,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n76,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n75,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n74,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n73,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n72,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n71,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n70,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n69,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n68,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n67,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n66,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n65,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n64,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n63,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n62,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n61,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n60,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n59,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n58,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n57,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n56,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n55,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n54,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n53,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n52,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n51,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n50,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n49,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n48,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n47,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n46,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n45,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n44,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n43,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n42,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n41,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n40,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n39,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n38,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n37,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n36,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n35,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n34,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n33,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n32,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n31,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n30,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n29,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n28,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n27,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n26,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n25,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n24,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n23,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n22,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n21,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n20,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n19,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n18,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n17,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n16,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n15,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n14,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n13,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n12,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n11,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n10,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n9,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n8,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n7,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n6,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n5,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n4,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n3,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n157,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n156,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n155,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n154,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n153,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n152,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n151,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n150,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n149,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n148,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n147,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n146,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n145,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n143,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n141,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n140,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n139,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n138,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n137,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n136,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n135,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n134,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n133,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n132,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n131,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n130,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n129,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n128,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n127,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n126,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n124,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n123,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n122,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n121,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n120,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n119,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n118,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n117,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n116,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n115,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n114,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n113,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n112,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n111,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n110,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n109,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n108,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n107,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n106,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n105,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n104,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n103,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n102,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n101,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n100,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n41,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n40,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n39,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n38,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n37,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n36,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n35,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n33,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n32,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n31,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n30,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n29,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n28,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n27,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n26,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n25,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n24,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n23,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n22,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n21,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n20,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n19,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n18,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n17,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n16,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n15,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n14,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n13,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n12,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n11,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n10,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n9,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n8,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n7,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n6,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n5,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n4,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n3,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_result_LE,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_N35,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_2_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_3_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_4_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_5_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_7_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_8_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_9_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_10_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_11_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_12_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_13_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_14_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_15_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_16_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_17_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_18_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_19_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_20_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_21_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_22_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_23_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_24_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_25_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_rst_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_rst_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_int_LE,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_2_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_3_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_4_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_5_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_7_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_8_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_9_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_10_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_11_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_12_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op2_int_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op1_int_6_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_1_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_18_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_19_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_20_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_21_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_22_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_23_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n10,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n9,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n8,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n7,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n6,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_SUM_14_,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_int_LE_FF_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_RST_FFX_1_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_RST_FFX_2_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_RST_FFX_2_Q,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_result_LE_FF_n1,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n152,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n151,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n150,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n149,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n148,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n147,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n146,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n145,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n144,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n143,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n142,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n141,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n140,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n139,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n138,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n137,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n136,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n135,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n134,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n133,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n132,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n131,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n130,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n129,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n128,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n127,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n126,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n125,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n124,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n123,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n122,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n121,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n120,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n119,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n118,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n117,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n116,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n115,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n114,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n113,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n112,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n111,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n110,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n109,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n108,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n107,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n106,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n105,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n104,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n103,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n102,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n101,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n100,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n99,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n98,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n97,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n96,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n95,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n94,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n93,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n92,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n91,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n90,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n89,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n88,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n87,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n86,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n85,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n84,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n83,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n82,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n81,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n74,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n72,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n181,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n180,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n179,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n178,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n177,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n176,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n175,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n174,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n173,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n172,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n171,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n170,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n169,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n168,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n120,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n119,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n118,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n117,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n116,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n115,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n114,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n113,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n112,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n111,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n110,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n109,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n108,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n107,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n106,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n105,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n104,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n103,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n102,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n101,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n100,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n99,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n98,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n97,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n95,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n94,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n93,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n92,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n91,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n90,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n89,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n88,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n87,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n86,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n85,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n83,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n82,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n81,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n80,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n79,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n78,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n77,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n76,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n75,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n74,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n73,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n72,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n71,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n70,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n69,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n68,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n67,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n66,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n65,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n64,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n63,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n62,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n61,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n60,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n59,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n58,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n57,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n56,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n55,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n54,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n53,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n52,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n51,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n50,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n49,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n48,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n47,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n46,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n45,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n44,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n43,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n42,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n41,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n40,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n39,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n38,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n37,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n36,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n35,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n34,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n33,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n32,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n31,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n30,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n29,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n28,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n27,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n26,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n25,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n24,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n23,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n22,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n21,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n20,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n19,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n18,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n17,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n16,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n15,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n14,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n13,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n12,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n11,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n10,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n9,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n8,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n7,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n6,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n5,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n4,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n3,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n2,
         extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n1,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n36,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n35,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n34,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n32,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n31,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n30,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n29,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n28,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n27,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n26,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n25,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n24,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n23,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n22,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n21,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n20,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n19,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n18,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n17,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n16,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n15,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n14,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n13,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n12,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n11,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n10,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n9,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n8,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n7,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n6,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n5,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n4,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n3,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n2,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n1,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n69,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n68,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n67,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n66,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n65,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n64,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n63,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n62,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n61,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n60,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n59,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n58,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n57,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n56,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n55,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n54,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n53,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n52,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n51,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n50,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n49,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n48,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n47,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n46,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n45,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n44,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n43,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n42,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n41,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n40,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n39,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n38,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n37,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n36,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n35,
         extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n92,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n91,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n90,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n89,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n88,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n87,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n86,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n85,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n84,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n83,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n82,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n81,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n80,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n79,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n77,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n76,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n75,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n74,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n73,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n72,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n71,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n70,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n69,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n68,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n67,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n66,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n65,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n64,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n63,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n62,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n61,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n60,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n59,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n58,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n57,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n56,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n55,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n54,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n53,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n52,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n51,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n50,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n49,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n48,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n47,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n46,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n45,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n44,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n43,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n40,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n1,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n78,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n41,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n39,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n38,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n37,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n36,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n35,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n34,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n33,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n32,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n31,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n30,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n29,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n28,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n27,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n26,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n25,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n24,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n23,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n22,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n21,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n20,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n19,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n18,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n17,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n16,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n15,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n14,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n13,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n12,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n11,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n10,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n9,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n8,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n7,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n6,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n5,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n4,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n3,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n2,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_0_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_1_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_2_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_3_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_4_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_5_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_6_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_7_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_8_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_9_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_10_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_11_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_12_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_13_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_14_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_15_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_16_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_17_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_18_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_19_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_n1,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_SUM_20_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n66,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n62,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n60,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n61,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n59,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n58,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n57,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n56,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n55,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n54,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n53,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n52,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n51,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n50,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n49,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n48,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n47,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n46,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n45,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n44,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n43,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n42,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n41,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n40,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n39,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n38,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n37,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n36,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n35,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n34,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n33,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n32,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n31,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n30,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n29,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n28,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n27,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n26,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n25,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n24,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n23,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n22,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n21,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n20,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n19,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n18,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n17,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n16,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n15,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n14,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n13,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n12,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n11,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n10,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n9,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n8,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n7,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n6,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n5,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n4,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n3,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n2,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n1,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n132,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n131,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n130,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n129,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n128,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n127,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n126,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n125,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n124,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n123,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n122,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n121,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n120,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n119,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n118,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n117,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n116,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n115,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n114,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n113,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n112,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n111,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n110,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n109,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n108,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n107,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n106,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n105,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n104,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n103,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n102,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n101,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n100,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n99,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n98,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n97,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n96,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n95,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n94,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n93,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n92,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n91,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n90,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n89,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n88,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n87,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n86,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n85,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n84,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n83,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n82,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n81,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n80,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n79,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n77,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n76,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n75,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n74,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n73,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n72,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n71,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n70,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n69,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n68,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n67,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n66,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n65,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n64,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n63,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n62,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n61,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n60,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n59,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n58,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n57,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n56,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n55,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n54,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n53,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n52,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n51,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n50,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n49,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n48,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n47,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n46,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n45,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n44,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n43,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n40,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n1,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_0_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_1_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_2_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_3_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_4_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_5_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_6_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_7_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_8_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_9_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_10_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_11_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_12_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_13_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_14_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_15_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_16_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_17_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_18_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_19_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_n1,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_SUM_20_,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n127,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n126,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n125,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n124,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n123,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n122,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n121,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n120,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n119,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n118,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n117,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n116,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n115,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n114,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n113,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n112,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n111,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n110,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n109,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n108,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n107,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n106,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n105,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n104,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n103,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n102,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n101,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n100,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n99,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n98,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n97,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n96,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n95,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n94,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n93,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n92,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n91,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n90,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n89,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n88,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n87,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n86,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n85,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n84,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n83,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n82,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n81,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n80,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n79,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n78,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n77,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n76,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n75,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n74,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n73,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n72,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n71,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n70,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n69,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n68,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n66,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n62,
         extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n60,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n26,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n25,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n12,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n11,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n10,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n9,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n8,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n7,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n6,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n5,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n2,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n1,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n4,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n3,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_N2,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_N0,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n28,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n27,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n26,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n25,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n12,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n11,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n10,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n9,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n8,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n7,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n6,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n5,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n2,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n1,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_N2,
         extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_N0,
         extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1,
         extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1,
         extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_n1,
         extimating_unit_Pixel_Retrieval_Unit_y_counter_n2,
         extimating_unit_Pixel_Retrieval_Unit_y_counter_n7,
         extimating_unit_Pixel_Retrieval_Unit_y_counter_n5,
         extimating_unit_Pixel_Retrieval_Unit_y_counter_n3,
         extimating_unit_Pixel_Retrieval_Unit_y_counter_n1,
         extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_n1,
         extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_n1,
         extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_n1,
         extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1,
         extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1,
         extimating_unit_extimator_CU_n31, extimating_unit_extimator_CU_n27,
         extimating_unit_extimator_CU_n23, extimating_unit_extimator_CU_n22,
         extimating_unit_extimator_CU_n21, extimating_unit_extimator_CU_n17,
         extimating_unit_extimator_CU_n15, extimating_unit_extimator_CU_n13,
         extimating_unit_extimator_CU_n12, extimating_unit_extimator_CU_n8,
         extimating_unit_extimator_CU_n7, extimating_unit_extimator_CU_n6,
         extimating_unit_extimator_CU_n5, extimating_unit_extimator_CU_n4,
         extimating_unit_extimator_CU_n3, extimating_unit_extimator_CU_n2,
         extimating_unit_extimator_CU_n1, extimating_unit_extimator_CU_n98,
         extimating_unit_extimator_CU_n97, extimating_unit_extimator_CU_n96,
         extimating_unit_extimator_CU_n95, extimating_unit_extimator_CU_n94,
         extimating_unit_extimator_CU_n93, extimating_unit_extimator_CU_n92,
         extimating_unit_extimator_CU_n91, extimating_unit_extimator_CU_n90,
         extimating_unit_extimator_CU_n89, extimating_unit_extimator_CU_n88,
         extimating_unit_extimator_CU_n87, extimating_unit_extimator_CU_n86,
         extimating_unit_extimator_CU_n85, extimating_unit_extimator_CU_n84,
         extimating_unit_extimator_CU_n83, extimating_unit_extimator_CU_n82,
         extimating_unit_extimator_CU_n81, extimating_unit_extimator_CU_n80,
         extimating_unit_extimator_CU_n79, extimating_unit_extimator_CU_n78,
         extimating_unit_extimator_CU_n77, extimating_unit_extimator_CU_n76,
         extimating_unit_extimator_CU_n75, extimating_unit_extimator_CU_n74,
         extimating_unit_extimator_CU_n73, extimating_unit_extimator_CU_n72,
         extimating_unit_extimator_CU_n71, extimating_unit_extimator_CU_n70,
         extimating_unit_extimator_CU_n69, extimating_unit_extimator_CU_n68,
         extimating_unit_extimator_CU_n67, extimating_unit_extimator_CU_n66,
         extimating_unit_extimator_CU_n65, extimating_unit_extimator_CU_n64,
         extimating_unit_extimator_CU_n63, extimating_unit_extimator_CU_n62,
         extimating_unit_extimator_CU_n61, extimating_unit_extimator_CU_n60,
         extimating_unit_extimator_CU_n59, extimating_unit_extimator_CU_n58,
         extimating_unit_extimator_CU_n57, extimating_unit_extimator_CU_n56,
         extimating_unit_extimator_CU_n55, extimating_unit_extimator_CU_n54,
         extimating_unit_extimator_CU_n53, extimating_unit_extimator_CU_n52,
         extimating_unit_extimator_CU_n51, extimating_unit_extimator_CU_n50,
         extimating_unit_extimator_CU_n49, extimating_unit_extimator_CU_n48,
         extimating_unit_extimator_CU_n47, extimating_unit_extimator_CU_n46,
         extimating_unit_extimator_CU_n45, extimating_unit_extimator_CU_n44,
         extimating_unit_extimator_CU_n43, extimating_unit_extimator_CU_n42,
         extimating_unit_extimator_CU_n41, extimating_unit_extimator_CU_n40,
         extimating_unit_extimator_CU_n39, extimating_unit_extimator_CU_n38,
         extimating_unit_extimator_CU_n37, extimating_unit_extimator_CU_n36,
         extimating_unit_extimator_CU_n35, extimating_unit_extimator_CU_n34,
         extimating_unit_extimator_CU_n33, extimating_unit_extimator_CU_n30,
         extimating_unit_extimator_CU_n29, extimating_unit_extimator_CU_n28,
         extimating_unit_extimator_CU_n25, extimating_unit_extimator_CU_n24,
         extimating_unit_extimator_CU_N183, extimating_unit_extimator_CU_N182,
         extimating_unit_extimator_CU_N181, extimating_unit_extimator_CU_N180,
         extimating_unit_extimator_CU_N179,
         extimating_unit_extimator_CU_CountTerm_OUT_int,
         extimating_unit_extimator_CU_Second_ready_int,
         extimating_unit_extimator_CU_last_cand_int,
         extimating_unit_extimator_CU_last_block_y_int,
         extimating_unit_extimator_CU_last_block_x_int,
         extimating_unit_extimator_CU_VALID_int,
         extimating_unit_extimator_CU_VALID_samp_n1,
         extimating_unit_extimator_CU_last_block_x_samp_n1,
         extimating_unit_extimator_CU_last_block_y_samp_n1,
         extimating_unit_extimator_CU_last_cand_samp_n1,
         extimating_unit_extimator_CU_Second_ready_samp_n1,
         extimating_unit_extimator_CU_CountTerm_OUT_samp_n1,
         extimating_unit_Ready_Handler_n4, extimating_unit_Ready_Handler_n2,
         extimating_unit_Ready_Handler_n1, extimating_unit_Ready_Handler_n9,
         extimating_unit_Ready_Handler_n8, extimating_unit_Ready_Handler_n7,
         extimating_unit_Ready_Handler_n6, extimating_unit_Ready_Handler_n5,
         extimating_unit_Ready_Handler_n3, extimating_unit_Ready_Handler_PS_0_,
         extimating_unit_Ready_Handler_PS_1_,
         extimating_unit_Ready_Handler_PS_2_, extimating_unit_CU_adapter_n14,
         extimating_unit_CU_adapter_n13, extimating_unit_CU_adapter_n12,
         extimating_unit_CU_adapter_n11, extimating_unit_CU_adapter_n10,
         extimating_unit_CU_adapter_n9, extimating_unit_CU_adapter_n6,
         extimating_unit_CU_adapter_n5, extimating_unit_CU_adapter_n4,
         extimating_unit_CU_adapter_n3, extimating_unit_CU_adapter_n2,
         extimating_unit_CU_adapter_n8, extimating_unit_CU_adapter_n7,
         extimating_unit_CU_adapter_n1,
         extimating_unit_CU_adapter_A3MVin_LE_samp,
         extimating_unit_CU_adapter_ADD3_MVin_LE_fRESET_half_delayed,
         extimating_unit_CU_adapter_MULT1_VALID_int_0_,
         extimating_unit_CU_adapter_MULT1_VALID_int_1_,
         extimating_unit_CU_adapter_idv_sel,
         extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_delay_1_n1,
         extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_delay_2_n1,
         extimating_unit_CU_adapter_inter_data_valid_FlFl_n1,
         extimating_unit_CU_adapter_MULT1_VALID_delay_1_n1,
         extimating_unit_CU_adapter_MULT1_VALID_delay_2_n1,
         extimating_unit_CU_adapter_ADD3_VALID_delay_1_n1,
         extimating_unit_CU_adapter_ADD3_VALID_delay_2_n1,
         extimating_unit_CU_adapter_ADD3_VALID_delay_3_n1,
         extimating_unit_CU_adapter_ADD3_VALID_delay_4_n1,
         extimating_unit_CU_adapter_ADD3_VALID_delay_5_n1,
         extimating_unit_CU_adapter_incrY_delay_1_n1,
         extimating_unit_CU_adapter_incrY_delay_2_n1,
         extimating_unit_CU_adapter_incrY_delay_3_n1,
         extimating_unit_CU_adapter_MEM_RE_delay_1_n1,
         extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_1_n1,
         extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_2_n1,
         extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_3_n1,
         extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_4_n1,
         extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_5_n1,
         extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_6_n1,
         extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_7_n1,
         extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_8_n1,
         extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_9_n1,
         extimating_unit_CU_adapter_ADD3_MVin_LE_register_n1,
         extimating_unit_CU_adapter_LE_ab_delay_1_n1,
         extimating_unit_CU_adapter_LE_ab_delay_2_n1,
         extimating_unit_CU_adapter_LE_ab_delay_3_n1,
         extimating_unit_CU_adapter_LE_ab_delay_4_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_1_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_2_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_3_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_4_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_5_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_6_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_7_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_8_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_9_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_10_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_11_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_12_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_13_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_14_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_15_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_16_n1,
         extimating_unit_CU_adapter_SAD_tmp_RST_delay_17_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_1_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_2_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_3_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_4_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_5_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_6_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_7_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_8_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_9_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_10_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_11_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_12_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_13_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_14_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_15_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_16_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_17_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_18_n1,
         extimating_unit_CU_adapter_Comp_EN_delay_19_n1,
         extimating_unit_Results_calculator_n217,
         extimating_unit_Results_calculator_n216,
         extimating_unit_Results_calculator_n215,
         extimating_unit_Results_calculator_n214,
         extimating_unit_Results_calculator_n213,
         extimating_unit_Results_calculator_n212,
         extimating_unit_Results_calculator_n211,
         extimating_unit_Results_calculator_n210,
         extimating_unit_Results_calculator_n209,
         extimating_unit_Results_calculator_n208,
         extimating_unit_Results_calculator_n207,
         extimating_unit_Results_calculator_n206,
         extimating_unit_Results_calculator_n205,
         extimating_unit_Results_calculator_n204,
         extimating_unit_Results_calculator_n203,
         extimating_unit_Results_calculator_n202,
         extimating_unit_Results_calculator_n201,
         extimating_unit_Results_calculator_n198,
         extimating_unit_Results_calculator_n199,
         extimating_unit_Results_calculator_n197,
         extimating_unit_Results_calculator_n196,
         extimating_unit_Results_calculator_n195,
         extimating_unit_Results_calculator_n194,
         extimating_unit_Results_calculator_n193,
         extimating_unit_Results_calculator_n192,
         extimating_unit_Results_calculator_n191,
         extimating_unit_Results_calculator_n190,
         extimating_unit_Results_calculator_n189,
         extimating_unit_Results_calculator_n188,
         extimating_unit_Results_calculator_n187,
         extimating_unit_Results_calculator_n186,
         extimating_unit_Results_calculator_n185,
         extimating_unit_Results_calculator_n184,
         extimating_unit_Results_calculator_n183,
         extimating_unit_Results_calculator_n182,
         extimating_unit_Results_calculator_n181,
         extimating_unit_Results_calculator_n180,
         extimating_unit_Results_calculator_n179,
         extimating_unit_Results_calculator_n178,
         extimating_unit_Results_calculator_n177,
         extimating_unit_Results_calculator_n176,
         extimating_unit_Results_calculator_n175,
         extimating_unit_Results_calculator_n174,
         extimating_unit_Results_calculator_n173,
         extimating_unit_Results_calculator_n172,
         extimating_unit_Results_calculator_n171,
         extimating_unit_Results_calculator_n170,
         extimating_unit_Results_calculator_n169,
         extimating_unit_Results_calculator_n168,
         extimating_unit_Results_calculator_n167,
         extimating_unit_Results_calculator_n166,
         extimating_unit_Results_calculator_n165,
         extimating_unit_Results_calculator_n164,
         extimating_unit_Results_calculator_n163,
         extimating_unit_Results_calculator_n162,
         extimating_unit_Results_calculator_n161,
         extimating_unit_Results_calculator_n160,
         extimating_unit_Results_calculator_n159,
         extimating_unit_Results_calculator_n158,
         extimating_unit_Results_calculator_n157,
         extimating_unit_Results_calculator_n156,
         extimating_unit_Results_calculator_n155,
         extimating_unit_Results_calculator_n154,
         extimating_unit_Results_calculator_n153,
         extimating_unit_Results_calculator_n152,
         extimating_unit_Results_calculator_n151,
         extimating_unit_Results_calculator_n150,
         extimating_unit_Results_calculator_n149,
         extimating_unit_Results_calculator_n148,
         extimating_unit_Results_calculator_n147,
         extimating_unit_Results_calculator_n146,
         extimating_unit_Results_calculator_n145,
         extimating_unit_Results_calculator_n144,
         extimating_unit_Results_calculator_n143,
         extimating_unit_Results_calculator_n142,
         extimating_unit_Results_calculator_n141,
         extimating_unit_Results_calculator_n140,
         extimating_unit_Results_calculator_n139,
         extimating_unit_Results_calculator_n138,
         extimating_unit_Results_calculator_n137,
         extimating_unit_Results_calculator_n136,
         extimating_unit_Results_calculator_n135,
         extimating_unit_Results_calculator_n134,
         extimating_unit_Results_calculator_n133,
         extimating_unit_Results_calculator_n132,
         extimating_unit_Results_calculator_n131,
         extimating_unit_Results_calculator_n130,
         extimating_unit_Results_calculator_n129,
         extimating_unit_Results_calculator_n128,
         extimating_unit_Results_calculator_n127,
         extimating_unit_Results_calculator_n126,
         extimating_unit_Results_calculator_n125,
         extimating_unit_Results_calculator_n124,
         extimating_unit_Results_calculator_n123,
         extimating_unit_Results_calculator_n122,
         extimating_unit_Results_calculator_n121,
         extimating_unit_Results_calculator_n120,
         extimating_unit_Results_calculator_n119,
         extimating_unit_Results_calculator_n118,
         extimating_unit_Results_calculator_n117,
         extimating_unit_Results_calculator_n116,
         extimating_unit_Results_calculator_n115,
         extimating_unit_Results_calculator_n114,
         extimating_unit_Results_calculator_n113,
         extimating_unit_Results_calculator_n112,
         extimating_unit_Results_calculator_n111,
         extimating_unit_Results_calculator_n110,
         extimating_unit_Results_calculator_n109,
         extimating_unit_Results_calculator_n108,
         extimating_unit_Results_calculator_n107,
         extimating_unit_Results_calculator_n106,
         extimating_unit_Results_calculator_n105,
         extimating_unit_Results_calculator_n104,
         extimating_unit_Results_calculator_n103,
         extimating_unit_Results_calculator_n102,
         extimating_unit_Results_calculator_n101,
         extimating_unit_Results_calculator_n100,
         extimating_unit_Results_calculator_n99,
         extimating_unit_Results_calculator_n98,
         extimating_unit_Results_calculator_n97,
         extimating_unit_Results_calculator_n96,
         extimating_unit_Results_calculator_n95,
         extimating_unit_Results_calculator_n94,
         extimating_unit_Results_calculator_n93,
         extimating_unit_Results_calculator_n92,
         extimating_unit_Results_calculator_n91,
         extimating_unit_Results_calculator_n90,
         extimating_unit_Results_calculator_n89,
         extimating_unit_Results_calculator_n88,
         extimating_unit_Results_calculator_n87,
         extimating_unit_Results_calculator_n86,
         extimating_unit_Results_calculator_n85,
         extimating_unit_Results_calculator_n84,
         extimating_unit_Results_calculator_n83,
         extimating_unit_Results_calculator_n82,
         extimating_unit_Results_calculator_n81,
         extimating_unit_Results_calculator_n80,
         extimating_unit_Results_calculator_n79,
         extimating_unit_Results_calculator_n78,
         extimating_unit_Results_calculator_n77,
         extimating_unit_Results_calculator_n76,
         extimating_unit_Results_calculator_n75,
         extimating_unit_Results_calculator_n74,
         extimating_unit_Results_calculator_n73,
         extimating_unit_Results_calculator_n72,
         extimating_unit_Results_calculator_n71,
         extimating_unit_Results_calculator_n70,
         extimating_unit_Results_calculator_n69,
         extimating_unit_Results_calculator_n68,
         extimating_unit_Results_calculator_n67,
         extimating_unit_Results_calculator_n66,
         extimating_unit_Results_calculator_n65,
         extimating_unit_Results_calculator_n64,
         extimating_unit_Results_calculator_n63,
         extimating_unit_Results_calculator_n62,
         extimating_unit_Results_calculator_n61,
         extimating_unit_Results_calculator_n60,
         extimating_unit_Results_calculator_n59,
         extimating_unit_Results_calculator_n58,
         extimating_unit_Results_calculator_n57,
         extimating_unit_Results_calculator_n56,
         extimating_unit_Results_calculator_n55,
         extimating_unit_Results_calculator_n54,
         extimating_unit_Results_calculator_n53,
         extimating_unit_Results_calculator_n52,
         extimating_unit_Results_calculator_n51,
         extimating_unit_Results_calculator_n50,
         extimating_unit_Results_calculator_n49,
         extimating_unit_Results_calculator_n48,
         extimating_unit_Results_calculator_n47,
         extimating_unit_Results_calculator_n46,
         extimating_unit_Results_calculator_n45,
         extimating_unit_Results_calculator_n44,
         extimating_unit_Results_calculator_n43,
         extimating_unit_Results_calculator_n42,
         extimating_unit_Results_calculator_n41,
         extimating_unit_Results_calculator_n40,
         extimating_unit_Results_calculator_n39,
         extimating_unit_Results_calculator_n38,
         extimating_unit_Results_calculator_n37,
         extimating_unit_Results_calculator_n36,
         extimating_unit_Results_calculator_n35,
         extimating_unit_Results_calculator_n34,
         extimating_unit_Results_calculator_n33,
         extimating_unit_Results_calculator_n32,
         extimating_unit_Results_calculator_n31,
         extimating_unit_Results_calculator_n30,
         extimating_unit_Results_calculator_n29,
         extimating_unit_Results_calculator_n28,
         extimating_unit_Results_calculator_n27,
         extimating_unit_Results_calculator_n26,
         extimating_unit_Results_calculator_n25,
         extimating_unit_Results_calculator_n24,
         extimating_unit_Results_calculator_n23,
         extimating_unit_Results_calculator_n22,
         extimating_unit_Results_calculator_n21,
         extimating_unit_Results_calculator_n20,
         extimating_unit_Results_calculator_n19,
         extimating_unit_Results_calculator_n18,
         extimating_unit_Results_calculator_n17,
         extimating_unit_Results_calculator_n16,
         extimating_unit_Results_calculator_n15,
         extimating_unit_Results_calculator_n14,
         extimating_unit_Results_calculator_n13,
         extimating_unit_Results_calculator_n12,
         extimating_unit_Results_calculator_n11,
         extimating_unit_Results_calculator_n10,
         extimating_unit_Results_calculator_n9,
         extimating_unit_Results_calculator_n8,
         extimating_unit_Results_calculator_n7,
         extimating_unit_Results_calculator_n6,
         extimating_unit_Results_calculator_n5,
         extimating_unit_Results_calculator_n4,
         extimating_unit_Results_calculator_n3,
         extimating_unit_Results_calculator_n2,
         extimating_unit_Results_calculator_n1,
         extimating_unit_Results_calculator_CurCand,
         extimating_unit_Results_calculator_Found_best,
         extimating_unit_Results_calculator_ltmin,
         extimating_unit_Results_calculator_CurSAD_tmp_0_,
         extimating_unit_Results_calculator_CurSAD_tmp_1_,
         extimating_unit_Results_calculator_CurSAD_tmp_2_,
         extimating_unit_Results_calculator_CurSAD_tmp_3_,
         extimating_unit_Results_calculator_CurSAD_tmp_4_,
         extimating_unit_Results_calculator_CurSAD_tmp_5_,
         extimating_unit_Results_calculator_CurSAD_tmp_6_,
         extimating_unit_Results_calculator_CurSAD_tmp_7_,
         extimating_unit_Results_calculator_CurSAD_tmp_8_,
         extimating_unit_Results_calculator_CurSAD_tmp_9_,
         extimating_unit_Results_calculator_CurSAD_tmp_10_,
         extimating_unit_Results_calculator_CurSAD_tmp_11_,
         extimating_unit_Results_calculator_CurSAD_tmp_12_,
         extimating_unit_Results_calculator_CurSAD_tmp_13_,
         extimating_unit_Results_calculator_CurSAD_tmp_14_,
         extimating_unit_Results_calculator_CurSAD_tmp_15_,
         extimating_unit_Results_calculator_CurSAD_tmp_16_,
         extimating_unit_Results_calculator_CurSAD_tmp_17_,
         extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n10,
         extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n9,
         extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n8,
         extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n7,
         extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n6,
         extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n5,
         extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n4,
         extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n3,
         extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n1,
         extimating_unit_Results_calculator_Pel_diff_reg_0_n1,
         extimating_unit_Results_calculator_Abs_X_0_n38,
         extimating_unit_Results_calculator_Abs_X_0_n29,
         extimating_unit_Results_calculator_Abs_X_0_n28,
         extimating_unit_Results_calculator_Abs_X_0_n27,
         extimating_unit_Results_calculator_Abs_X_0_n26,
         extimating_unit_Results_calculator_Abs_X_0_n25,
         extimating_unit_Results_calculator_Abs_X_0_n24,
         extimating_unit_Results_calculator_Abs_X_0_n23,
         extimating_unit_Results_calculator_Abs_X_0_n22,
         extimating_unit_Results_calculator_Abs_X_0_n13,
         extimating_unit_Results_calculator_Abs_X_0_n12,
         extimating_unit_Results_calculator_Abs_X_0_n11,
         extimating_unit_Results_calculator_Abs_X_0_n10,
         extimating_unit_Results_calculator_Abs_X_0_n9,
         extimating_unit_Results_calculator_Abs_X_0_n8,
         extimating_unit_Results_calculator_Abs_X_0_n7,
         extimating_unit_Results_calculator_Abs_X_0_n6,
         extimating_unit_Results_calculator_Abs_X_0_n5,
         extimating_unit_Results_calculator_Abs_X_0_n4,
         extimating_unit_Results_calculator_Abs_X_0_n3,
         extimating_unit_Results_calculator_Abs_X_0_n2,
         extimating_unit_Results_calculator_Abs_X_0_n1,
         extimating_unit_Results_calculator_Abs_X_0_n21,
         extimating_unit_Results_calculator_Abs_X_0_n20,
         extimating_unit_Results_calculator_Abs_X_0_n19,
         extimating_unit_Results_calculator_Abs_X_0_n18,
         extimating_unit_Results_calculator_Abs_X_0_n17,
         extimating_unit_Results_calculator_Abs_X_0_n16,
         extimating_unit_Results_calculator_Abs_X_0_n15,
         extimating_unit_Results_calculator_Abs_X_0_n14,
         extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_n1,
         extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n10,
         extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n9,
         extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n8,
         extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n7,
         extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n6,
         extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n5,
         extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n4,
         extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n3,
         extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n1,
         extimating_unit_Results_calculator_Pel_diff_reg_1_n1,
         extimating_unit_Results_calculator_Abs_X_1_n46,
         extimating_unit_Results_calculator_Abs_X_1_n45,
         extimating_unit_Results_calculator_Abs_X_1_n44,
         extimating_unit_Results_calculator_Abs_X_1_n43,
         extimating_unit_Results_calculator_Abs_X_1_n42,
         extimating_unit_Results_calculator_Abs_X_1_n41,
         extimating_unit_Results_calculator_Abs_X_1_n40,
         extimating_unit_Results_calculator_Abs_X_1_n39,
         extimating_unit_Results_calculator_Abs_X_1_n38,
         extimating_unit_Results_calculator_Abs_X_1_n29,
         extimating_unit_Results_calculator_Abs_X_1_n28,
         extimating_unit_Results_calculator_Abs_X_1_n27,
         extimating_unit_Results_calculator_Abs_X_1_n26,
         extimating_unit_Results_calculator_Abs_X_1_n25,
         extimating_unit_Results_calculator_Abs_X_1_n24,
         extimating_unit_Results_calculator_Abs_X_1_n23,
         extimating_unit_Results_calculator_Abs_X_1_n22,
         extimating_unit_Results_calculator_Abs_X_1_n13,
         extimating_unit_Results_calculator_Abs_X_1_n12,
         extimating_unit_Results_calculator_Abs_X_1_n11,
         extimating_unit_Results_calculator_Abs_X_1_n10,
         extimating_unit_Results_calculator_Abs_X_1_n9,
         extimating_unit_Results_calculator_Abs_X_1_n8,
         extimating_unit_Results_calculator_Abs_X_1_n7,
         extimating_unit_Results_calculator_Abs_X_1_n6,
         extimating_unit_Results_calculator_Abs_X_1_n5,
         extimating_unit_Results_calculator_Abs_X_1_n4,
         extimating_unit_Results_calculator_Abs_X_1_n3,
         extimating_unit_Results_calculator_Abs_X_1_n2,
         extimating_unit_Results_calculator_Abs_X_1_n1,
         extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_n1,
         extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n10,
         extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n9,
         extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n8,
         extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n7,
         extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n6,
         extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n5,
         extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n4,
         extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n3,
         extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n1,
         extimating_unit_Results_calculator_Pel_diff_reg_2_n1,
         extimating_unit_Results_calculator_Abs_X_2_n46,
         extimating_unit_Results_calculator_Abs_X_2_n45,
         extimating_unit_Results_calculator_Abs_X_2_n44,
         extimating_unit_Results_calculator_Abs_X_2_n43,
         extimating_unit_Results_calculator_Abs_X_2_n42,
         extimating_unit_Results_calculator_Abs_X_2_n41,
         extimating_unit_Results_calculator_Abs_X_2_n40,
         extimating_unit_Results_calculator_Abs_X_2_n39,
         extimating_unit_Results_calculator_Abs_X_2_n38,
         extimating_unit_Results_calculator_Abs_X_2_n29,
         extimating_unit_Results_calculator_Abs_X_2_n28,
         extimating_unit_Results_calculator_Abs_X_2_n27,
         extimating_unit_Results_calculator_Abs_X_2_n26,
         extimating_unit_Results_calculator_Abs_X_2_n25,
         extimating_unit_Results_calculator_Abs_X_2_n24,
         extimating_unit_Results_calculator_Abs_X_2_n23,
         extimating_unit_Results_calculator_Abs_X_2_n22,
         extimating_unit_Results_calculator_Abs_X_2_n13,
         extimating_unit_Results_calculator_Abs_X_2_n12,
         extimating_unit_Results_calculator_Abs_X_2_n11,
         extimating_unit_Results_calculator_Abs_X_2_n10,
         extimating_unit_Results_calculator_Abs_X_2_n9,
         extimating_unit_Results_calculator_Abs_X_2_n8,
         extimating_unit_Results_calculator_Abs_X_2_n7,
         extimating_unit_Results_calculator_Abs_X_2_n6,
         extimating_unit_Results_calculator_Abs_X_2_n5,
         extimating_unit_Results_calculator_Abs_X_2_n4,
         extimating_unit_Results_calculator_Abs_X_2_n3,
         extimating_unit_Results_calculator_Abs_X_2_n2,
         extimating_unit_Results_calculator_Abs_X_2_n1,
         extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_n1,
         extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n10,
         extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n9,
         extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n8,
         extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n7,
         extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n6,
         extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n5,
         extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n4,
         extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n3,
         extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n1,
         extimating_unit_Results_calculator_Pel_diff_reg_3_n1,
         extimating_unit_Results_calculator_Abs_X_3_n46,
         extimating_unit_Results_calculator_Abs_X_3_n45,
         extimating_unit_Results_calculator_Abs_X_3_n44,
         extimating_unit_Results_calculator_Abs_X_3_n43,
         extimating_unit_Results_calculator_Abs_X_3_n42,
         extimating_unit_Results_calculator_Abs_X_3_n41,
         extimating_unit_Results_calculator_Abs_X_3_n40,
         extimating_unit_Results_calculator_Abs_X_3_n39,
         extimating_unit_Results_calculator_Abs_X_3_n38,
         extimating_unit_Results_calculator_Abs_X_3_n29,
         extimating_unit_Results_calculator_Abs_X_3_n28,
         extimating_unit_Results_calculator_Abs_X_3_n27,
         extimating_unit_Results_calculator_Abs_X_3_n26,
         extimating_unit_Results_calculator_Abs_X_3_n25,
         extimating_unit_Results_calculator_Abs_X_3_n24,
         extimating_unit_Results_calculator_Abs_X_3_n23,
         extimating_unit_Results_calculator_Abs_X_3_n22,
         extimating_unit_Results_calculator_Abs_X_3_n13,
         extimating_unit_Results_calculator_Abs_X_3_n12,
         extimating_unit_Results_calculator_Abs_X_3_n11,
         extimating_unit_Results_calculator_Abs_X_3_n10,
         extimating_unit_Results_calculator_Abs_X_3_n9,
         extimating_unit_Results_calculator_Abs_X_3_n8,
         extimating_unit_Results_calculator_Abs_X_3_n7,
         extimating_unit_Results_calculator_Abs_X_3_n6,
         extimating_unit_Results_calculator_Abs_X_3_n5,
         extimating_unit_Results_calculator_Abs_X_3_n4,
         extimating_unit_Results_calculator_Abs_X_3_n3,
         extimating_unit_Results_calculator_Abs_X_3_n2,
         extimating_unit_Results_calculator_Abs_X_3_n1,
         extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_n1,
         extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_n1,
         extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_n1,
         extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_n1,
         extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_n1,
         extimating_unit_Results_calculator_PelAdd_stage2_add_23_n1,
         extimating_unit_Results_calculator_CurRowSAD_reg_n1,
         extimating_unit_Results_calculator_SAD_tmp_reg_n19,
         extimating_unit_Results_calculator_SAD_tmp_reg_n18,
         extimating_unit_Results_calculator_SAD_tmp_reg_n17,
         extimating_unit_Results_calculator_SAD_tmp_reg_n16,
         extimating_unit_Results_calculator_SAD_tmp_reg_n15,
         extimating_unit_Results_calculator_SAD_tmp_reg_n14,
         extimating_unit_Results_calculator_SAD_tmp_reg_n13,
         extimating_unit_Results_calculator_SAD_tmp_reg_n12,
         extimating_unit_Results_calculator_SAD_tmp_reg_n11,
         extimating_unit_Results_calculator_SAD_tmp_reg_n10,
         extimating_unit_Results_calculator_SAD_tmp_reg_n9,
         extimating_unit_Results_calculator_SAD_tmp_reg_n8,
         extimating_unit_Results_calculator_SAD_tmp_reg_n7,
         extimating_unit_Results_calculator_SAD_tmp_reg_n6,
         extimating_unit_Results_calculator_SAD_tmp_reg_n5,
         extimating_unit_Results_calculator_SAD_tmp_reg_n4,
         extimating_unit_Results_calculator_SAD_tmp_reg_n3,
         extimating_unit_Results_calculator_SAD_tmp_reg_n2,
         extimating_unit_Results_calculator_SAD_tmp_reg_n1,
         extimating_unit_Results_calculator_CurSAD_reg_n1,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n197,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n196,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n195,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n194,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n193,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n192,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n191,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n190,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n189,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n188,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n187,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n186,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n185,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n184,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n183,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n182,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n181,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n180,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n179,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n178,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n177,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n176,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n175,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n174,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n173,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n172,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n171,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n170,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n169,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n168,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n167,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n166,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n165,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n164,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n163,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n162,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n161,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n160,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n159,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n158,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n157,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n156,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n155,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n154,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n153,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n152,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n151,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n150,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n149,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n148,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n147,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n146,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n145,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n144,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n143,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n142,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n141,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n140,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n139,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n138,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n137,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n136,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n135,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n134,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n133,
         extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n132,
         extimating_unit_Results_calculator_SAD_min_register_n58,
         extimating_unit_Results_calculator_SAD_min_register_n57,
         extimating_unit_Results_calculator_SAD_min_register_n56,
         extimating_unit_Results_calculator_SAD_min_register_n54,
         extimating_unit_Results_calculator_SAD_min_register_n55,
         extimating_unit_Results_calculator_SAD_min_register_n53,
         extimating_unit_Results_calculator_SAD_min_register_n52,
         extimating_unit_Results_calculator_SAD_min_register_n51,
         extimating_unit_Results_calculator_SAD_min_register_n50,
         extimating_unit_Results_calculator_SAD_min_register_n49,
         extimating_unit_Results_calculator_SAD_min_register_n48,
         extimating_unit_Results_calculator_SAD_min_register_n47,
         extimating_unit_Results_calculator_SAD_min_register_n46,
         extimating_unit_Results_calculator_SAD_min_register_n45,
         extimating_unit_Results_calculator_SAD_min_register_n44,
         extimating_unit_Results_calculator_SAD_min_register_n43,
         extimating_unit_Results_calculator_SAD_min_register_n42,
         extimating_unit_Results_calculator_SAD_min_register_n41,
         extimating_unit_Results_calculator_SAD_min_register_n40,
         extimating_unit_Results_calculator_SAD_min_register_n39,
         extimating_unit_Results_calculator_SAD_min_register_n38,
         extimating_unit_Results_calculator_SAD_min_register_n37,
         extimating_unit_Results_calculator_SAD_min_register_n36,
         extimating_unit_Results_calculator_SAD_min_register_n35,
         extimating_unit_Results_calculator_SAD_min_register_n34,
         extimating_unit_Results_calculator_SAD_min_register_n33,
         extimating_unit_Results_calculator_SAD_min_register_n32,
         extimating_unit_Results_calculator_SAD_min_register_n31,
         extimating_unit_Results_calculator_SAD_min_register_n30,
         extimating_unit_Results_calculator_SAD_min_register_n29,
         extimating_unit_Results_calculator_SAD_min_register_n28,
         extimating_unit_Results_calculator_SAD_min_register_n27,
         extimating_unit_Results_calculator_SAD_min_register_n26,
         extimating_unit_Results_calculator_SAD_min_register_n25,
         extimating_unit_Results_calculator_SAD_min_register_n24,
         extimating_unit_Results_calculator_SAD_min_register_n23,
         extimating_unit_Results_calculator_SAD_min_register_n22,
         extimating_unit_Results_calculator_SAD_min_register_n21,
         extimating_unit_Results_calculator_SAD_min_register_n20,
         extimating_unit_Results_calculator_SAD_min_register_n19,
         extimating_unit_Results_calculator_SAD_min_register_n18,
         extimating_unit_Results_calculator_SAD_min_register_n17,
         extimating_unit_Results_calculator_SAD_min_register_n16,
         extimating_unit_Results_calculator_SAD_min_register_n15,
         extimating_unit_Results_calculator_SAD_min_register_n14,
         extimating_unit_Results_calculator_SAD_min_register_n13,
         extimating_unit_Results_calculator_SAD_min_register_n12,
         extimating_unit_Results_calculator_SAD_min_register_n11,
         extimating_unit_Results_calculator_SAD_min_register_n10,
         extimating_unit_Results_calculator_SAD_min_register_n9,
         extimating_unit_Results_calculator_SAD_min_register_n8,
         extimating_unit_Results_calculator_SAD_min_register_n7,
         extimating_unit_Results_calculator_SAD_min_register_n6,
         extimating_unit_Results_calculator_SAD_min_register_n5,
         extimating_unit_Results_calculator_SAD_min_register_n4,
         extimating_unit_Results_calculator_SAD_min_register_n3,
         extimating_unit_Results_calculator_SAD_min_register_n2,
         extimating_unit_Results_calculator_SAD_min_register_n1,
         extimating_unit_Results_calculator_CurCand_counter_n1,
         extimating_unit_Results_calculator_CurCand_counter_n2,
         extimating_unit_Results_calculator_BestCand_register_n3,
         extimating_unit_Results_calculator_BestCand_register_n4,
         extimating_unit_Results_calculator_BestCand_register_n2,
         extimating_unit_Results_calculator_BestCand_register_n1,
         extimating_unit_Results_calculator_Terminal_counter_n7,
         extimating_unit_Results_calculator_Terminal_counter_n18,
         extimating_unit_Results_calculator_Terminal_counter_n16,
         extimating_unit_Results_calculator_Terminal_counter_n15,
         extimating_unit_Results_calculator_Terminal_counter_n14,
         extimating_unit_Results_calculator_Terminal_counter_n13,
         extimating_unit_Results_calculator_Terminal_counter_n11,
         extimating_unit_Results_calculator_Terminal_counter_n10,
         extimating_unit_Results_calculator_Terminal_counter_n9,
         extimating_unit_Results_calculator_Terminal_counter_n8,
         extimating_unit_Results_calculator_Terminal_counter_n6,
         extimating_unit_Results_calculator_Terminal_counter_n5,
         extimating_unit_Results_calculator_Terminal_counter_n4,
         extimating_unit_Results_calculator_Terminal_counter_n3,
         extimating_unit_Results_calculator_Terminal_counter_n2,
         extimating_unit_Results_calculator_Terminal_counter_n1,
         extimating_unit_Results_calculator_Terminal_counter_N6,
         extimating_unit_Results_calculator_Terminal_counter_N5,
         extimating_unit_Results_calculator_Terminal_counter_N4,
         extimating_unit_Results_calculator_Terminal_counter_N3,
         extimating_unit_Results_calculator_Terminal_counter_N2,
         extimating_unit_Results_calculator_Terminal_counter_count_0_,
         extimating_unit_Results_calculator_Terminal_counter_count_1_,
         extimating_unit_Results_calculator_Terminal_counter_count_2_,
         extimating_unit_Results_calculator_Terminal_counter_count_3_,
         extimating_unit_Results_calculator_Terminal_counter_count_4_,
         extimating_unit_Results_calculator_Candidate_counter_n3,
         extimating_unit_Results_calculator_Candidate_counter_n1,
         extimating_unit_Results_calculator_add_85_n17,
         extimating_unit_Results_calculator_add_85_n7,
         extimating_unit_Results_calculator_add_85_n6,
         extimating_unit_Results_calculator_add_85_n5,
         extimating_unit_Results_calculator_add_85_n4,
         extimating_unit_Results_calculator_add_85_n3,
         extimating_unit_Results_calculator_add_85_n2,
         extimating_unit_Results_calculator_add_85_n1,
         extimating_unit_Results_calculator_add_85_carry_2_,
         extimating_unit_Results_calculator_add_85_carry_3_,
         extimating_unit_Results_calculator_add_85_carry_4_,
         extimating_unit_Results_calculator_add_85_carry_5_,
         extimating_unit_Results_calculator_add_85_carry_6_,
         extimating_unit_Results_calculator_add_85_carry_7_,
         extimating_unit_Results_calculator_add_85_carry_8_,
         extimating_unit_Results_calculator_add_85_carry_9_,
         extimating_unit_Results_calculator_add_85_carry_10_;
  wire   [2:0] constructing_unit_Control_Unit_NS;
  wire   [27:0] constructing_unit_Datapath_D_min;
  wire   [27:0] constructing_unit_Datapath_D_Cur_tmp;
  wire   [27:0] constructing_unit_Datapath_D_sq;
  wire   [26:0] constructing_unit_Datapath_D_v_sq;
  wire   [26:0] constructing_unit_Datapath_D_h_sq;
  wire   [2:0] constructing_unit_Datapath_UA_flag;
  wire   [26:0] constructing_unit_Datapath_D_v_sq_tmp;
  wire   [14:0] constructing_unit_Datapath_D_v_tmp;
  wire   [25:0] constructing_unit_Datapath_MV2_int_v_ext;
  wire   [29:0] constructing_unit_Datapath_MV2p_int_v;
  wire   [24:0] constructing_unit_Datapath_MV0_int_v_ext;
  wire   [27:0] constructing_unit_Datapath_diff_mult_h_int;
  wire   [59:0] constructing_unit_Datapath_mv1h_mv0h_int;
  wire   [26:0] constructing_unit_Datapath_D_h_sq_tmp;
  wire   [14:0] constructing_unit_Datapath_D_h_tmp;
  wire   [25:0] constructing_unit_Datapath_MV2_int_h_ext;
  wire   [29:0] constructing_unit_Datapath_MV2p_int_h;
  wire   [24:0] constructing_unit_Datapath_MV0_int_h_ext;
  wire   [27:0] constructing_unit_Datapath_diff_mult_v_int;
  wire   [1:0] constructing_unit_Datapath_CU_w_int;
  wire   [1:0] constructing_unit_Datapath_CU_h_int;
  wire   [59:0] constructing_unit_Datapath_mv1v_mv0v_int;
  wire   [11:1] constructing_unit_Datapath_L_sub1_sub_19_carry;
  wire   [1:0] constructing_unit_Datapath_hOw_cmd_RSH_out;
  wire   [1:0] constructing_unit_Datapath_hOw_RSH_in;
  wire   [2:1] constructing_unit_Datapath_hOw_shift_dir_int;
  wire   [13:0] constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L;
  wire   [12:0] constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L;
  wire   [13:0] constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext;
  wire   [11:0] constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R;
  wire   [14:1] constructing_unit_Datapath_L_sub2_sub_19_carry;
  wire   [14:1] constructing_unit_Datapath_L_subD_sub_19_carry;
  wire   [11:1] constructing_unit_Datapath_R_sub1_sub_19_carry;
  wire   [13:0] constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L;
  wire   [12:0] constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L;
  wire   [13:0] constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext;
  wire   [11:0] constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R;
  wire   [14:2] constructing_unit_Datapath_R_sum_add_19_carry;
  wire   [14:1] constructing_unit_Datapath_R_subD_sub_19_carry;
  wire   [27:2] constructing_unit_Datapath_D_adder_add_19_carry;
  wire   [1:0] extimating_unit_RF_Addr_CU_int;
  wire   [21:0] extimating_unit_MV2_out_int;
  wire   [21:0] extimating_unit_MV1_out_int;
  wire   [21:0] extimating_unit_MV0_out_int;
  wire   [12:0] extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp;
  wire   [12:0] extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp;
  wire   [11:0] extimating_unit_Pixel_Retrieval_Unit_MVr_h;
  wire   [11:0] extimating_unit_Pixel_Retrieval_Unit_MVr_v;
  wire   [11:0] extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp;
  wire   [11:0] extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp;
  wire   [19:0] extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h;
  wire   [19:0] extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v;
  wire   [21:0] extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext;
  wire   [17:0] extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3;
  wire   [17:0] extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2;
  wire   [17:0] extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1;
  wire   [17:0] extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0;
  wire   [47:0] extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp;
  wire   [11:1] extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv;
  wire   [47:0] extimating_unit_Pixel_Retrieval_Unit_R_SH2_out;
  wire   [7:0] extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp;
  wire   [47:0] extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp;
  wire   [47:0] extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp;
  wire  
         [1:0] extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_block_num
;
  wire  
         [1:0] extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_block_num
;
  wire   [11:1] extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry;
  wire   [11:1] extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry;
  wire   [11:1] extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry;
  wire   [11:1] extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry;
  wire   [11:0] extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int;
  wire   [11:0] extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int;
  wire   [11:0] extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int;
  wire   [11:0] extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int;
  wire   [13:0] extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1;
  wire   [13:0] extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int;
  wire  
         [13:2] extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry
;
  wire   [13:0] extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1;
  wire   [13:0] extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int;
  wire  
         [13:2] extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry
;
  wire   [13:0] extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1;
  wire   [13:0] extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int;
  wire  
         [13:2] extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry
;
  wire   [13:0] extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1;
  wire   [13:0] extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int;
  wire  
         [13:2] extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry
;
  wire   [19:0] extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp;
  wire  
         [19:2] extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry
;
  wire   [19:0] extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp;
  wire  
         [19:2] extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry
;
  wire  
         [12:2] extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry
;
  wire  
         [12:2] extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry
;
  wire   [11:2] extimating_unit_Pixel_Retrieval_Unit_add_140_carry;
  wire   [2:1] extimating_unit_Ready_Handler_NS;
  wire   [18:1] extimating_unit_CU_adapter_Comp_EN_int;
  wire   [16:1] extimating_unit_CU_adapter_SAD_tmp_RST_int;
  wire   [3:1] extimating_unit_CU_adapter_LE_ab_int;
  wire   [9:1] extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int;
  wire   [2:1] extimating_unit_CU_adapter_incrY_int;
  wire   [4:1] extimating_unit_CU_adapter_ADD3_VALID_int;
  wire   [2:1] extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_int;
  wire   [17:0] extimating_unit_Results_calculator_SAD_min;
  wire   [17:0] extimating_unit_Results_calculator_SAD_tmp;
  wire   [9:0] extimating_unit_Results_calculator_CurRowSAD;
  wire   [9:0] extimating_unit_Results_calculator_PelAdd_out;
  wire   [17:0] extimating_unit_Results_calculator_PelAdd_stage1_out_samp;
  wire   [17:0] extimating_unit_Results_calculator_PelAdd_stage1_out;
  wire   [31:0] extimating_unit_Results_calculator_ABs_Pel_diff_samp;
  wire   [31:0] extimating_unit_Results_calculator_Abs_Pel_diff;
  wire   [35:0] extimating_unit_Results_calculator_Pel_diff_samp;
  wire   [35:0] extimating_unit_Results_calculator_Pel_diff;
  wire   [8:1] extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry;
  wire   [8:1] extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry;
  wire   [8:1] extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry;
  wire   [8:1] extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry;
  wire  
         [7:2] extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_carry
;
  wire  
         [7:2] extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_carry
;
  wire   [8:2] extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry;
  wire  
         [2:4] extimating_unit_Results_calculator_Terminal_counter_add_23_carry
;
  assign Comp_EN = eComp_EN;
  assign CandCount_CE = ADD3_MVin_LE_nSET;
  assign RF_in_RE = 1'b1;

  INV_X1 U135 ( .A(n177), .ZN(n145) );
  INV_X1 U136 ( .A(n176), .ZN(n144) );
  INV_X1 U137 ( .A(n176), .ZN(n143) );
  INV_X1 U138 ( .A(n176), .ZN(n142) );
  INV_X1 U139 ( .A(n177), .ZN(n146) );
  BUF_X1 U140 ( .A(n140), .Z(n139) );
  BUF_X1 U141 ( .A(n140), .Z(n137) );
  BUF_X1 U142 ( .A(n140), .Z(n138) );
  BUF_X1 U143 ( .A(n141), .Z(n136) );
  BUF_X1 U144 ( .A(n141), .Z(n135) );
  INV_X1 U145 ( .A(n100), .ZN(n199) );
  AOI22_X1 U146 ( .A1(MVP1[11]), .A2(n144), .B1(eMV1_in[11]), .B2(n159), .ZN(
        n100) );
  INV_X1 U147 ( .A(n98), .ZN(n198) );
  AOI22_X1 U148 ( .A1(MVP1[12]), .A2(n144), .B1(eMV1_in[12]), .B2(n158), .ZN(
        n98) );
  INV_X1 U149 ( .A(n99), .ZN(n189) );
  AOI22_X1 U150 ( .A1(MVP1[21]), .A2(n144), .B1(eMV1_in[21]), .B2(n158), .ZN(
        n99) );
  INV_X1 U151 ( .A(n111), .ZN(n232) );
  AOI22_X1 U152 ( .A1(MVP1[0]), .A2(n143), .B1(eMV1_in[0]), .B2(n164), .ZN(
        n111) );
  INV_X1 U153 ( .A(n109), .ZN(n231) );
  AOI22_X1 U154 ( .A1(MVP1[1]), .A2(n144), .B1(eMV1_in[1]), .B2(n163), .ZN(
        n109) );
  INV_X1 U155 ( .A(n108), .ZN(n230) );
  AOI22_X1 U156 ( .A1(MVP1[2]), .A2(n144), .B1(eMV1_in[2]), .B2(n163), .ZN(
        n108) );
  INV_X1 U157 ( .A(n107), .ZN(n229) );
  AOI22_X1 U158 ( .A1(MVP1[3]), .A2(n144), .B1(eMV1_in[3]), .B2(n162), .ZN(
        n107) );
  INV_X1 U159 ( .A(n106), .ZN(n228) );
  AOI22_X1 U160 ( .A1(MVP1[4]), .A2(n144), .B1(eMV1_in[4]), .B2(n162), .ZN(
        n106) );
  INV_X1 U161 ( .A(n105), .ZN(n227) );
  AOI22_X1 U162 ( .A1(MVP1[5]), .A2(n144), .B1(eMV1_in[5]), .B2(n161), .ZN(
        n105) );
  INV_X1 U163 ( .A(n104), .ZN(n226) );
  AOI22_X1 U164 ( .A1(MVP1[6]), .A2(n144), .B1(eMV1_in[6]), .B2(n161), .ZN(
        n104) );
  INV_X1 U165 ( .A(n103), .ZN(n225) );
  AOI22_X1 U166 ( .A1(MVP1[7]), .A2(n144), .B1(eMV1_in[7]), .B2(n160), .ZN(
        n103) );
  INV_X1 U167 ( .A(n102), .ZN(n224) );
  AOI22_X1 U168 ( .A1(MVP1[8]), .A2(n144), .B1(eMV1_in[8]), .B2(n160), .ZN(
        n102) );
  INV_X1 U169 ( .A(n101), .ZN(n223) );
  AOI22_X1 U170 ( .A1(MVP1[9]), .A2(n144), .B1(eMV1_in[9]), .B2(n159), .ZN(
        n101) );
  INV_X1 U171 ( .A(n110), .ZN(n222) );
  AOI22_X1 U172 ( .A1(MVP1[10]), .A2(n143), .B1(eMV1_in[10]), .B2(n164), .ZN(
        n110) );
  INV_X1 U173 ( .A(n122), .ZN(n188) );
  AOI22_X1 U174 ( .A1(MVP0[11]), .A2(n142), .B1(eMV0_in[11]), .B2(n170), .ZN(
        n122) );
  INV_X1 U175 ( .A(n120), .ZN(n187) );
  AOI22_X1 U176 ( .A1(MVP0[12]), .A2(n143), .B1(eMV0_in[12]), .B2(n169), .ZN(
        n120) );
  INV_X1 U177 ( .A(n119), .ZN(n186) );
  AOI22_X1 U178 ( .A1(MVP0[13]), .A2(n143), .B1(eMV0_in[13]), .B2(n168), .ZN(
        n119) );
  INV_X1 U179 ( .A(n118), .ZN(n185) );
  AOI22_X1 U180 ( .A1(MVP0[14]), .A2(n143), .B1(eMV0_in[14]), .B2(n168), .ZN(
        n118) );
  INV_X1 U181 ( .A(n117), .ZN(n184) );
  AOI22_X1 U182 ( .A1(MVP0[15]), .A2(n143), .B1(eMV0_in[15]), .B2(n167), .ZN(
        n117) );
  INV_X1 U183 ( .A(n116), .ZN(n183) );
  AOI22_X1 U184 ( .A1(MVP0[16]), .A2(n143), .B1(eMV0_in[16]), .B2(n167), .ZN(
        n116) );
  INV_X1 U185 ( .A(n115), .ZN(n182) );
  AOI22_X1 U186 ( .A1(MVP0[17]), .A2(n143), .B1(eMV0_in[17]), .B2(n166), .ZN(
        n115) );
  INV_X1 U187 ( .A(n114), .ZN(n181) );
  AOI22_X1 U188 ( .A1(MVP0[18]), .A2(n143), .B1(eMV0_in[18]), .B2(n166), .ZN(
        n114) );
  INV_X1 U189 ( .A(n113), .ZN(n180) );
  AOI22_X1 U190 ( .A1(MVP0[19]), .A2(n143), .B1(eMV0_in[19]), .B2(n165), .ZN(
        n113) );
  INV_X1 U191 ( .A(n112), .ZN(n179) );
  AOI22_X1 U192 ( .A1(MVP0[20]), .A2(n143), .B1(eMV0_in[20]), .B2(n165), .ZN(
        n112) );
  INV_X1 U193 ( .A(n121), .ZN(n178) );
  AOI22_X1 U194 ( .A1(MVP0[21]), .A2(n143), .B1(eMV0_in[21]), .B2(n169), .ZN(
        n121) );
  INV_X1 U195 ( .A(n133), .ZN(n221) );
  AOI22_X1 U196 ( .A1(MVP0[0]), .A2(n142), .B1(eMV0_in[0]), .B2(n175), .ZN(
        n133) );
  INV_X1 U197 ( .A(n131), .ZN(n220) );
  AOI22_X1 U198 ( .A1(MVP0[1]), .A2(n142), .B1(eMV0_in[1]), .B2(n174), .ZN(
        n131) );
  INV_X1 U199 ( .A(n130), .ZN(n219) );
  AOI22_X1 U200 ( .A1(MVP0[2]), .A2(n142), .B1(eMV0_in[2]), .B2(n174), .ZN(
        n130) );
  INV_X1 U201 ( .A(n129), .ZN(n218) );
  AOI22_X1 U202 ( .A1(MVP0[3]), .A2(n142), .B1(eMV0_in[3]), .B2(n173), .ZN(
        n129) );
  INV_X1 U203 ( .A(n128), .ZN(n217) );
  AOI22_X1 U204 ( .A1(MVP0[4]), .A2(n142), .B1(eMV0_in[4]), .B2(n173), .ZN(
        n128) );
  INV_X1 U205 ( .A(n127), .ZN(n216) );
  AOI22_X1 U206 ( .A1(MVP0[5]), .A2(n142), .B1(eMV0_in[5]), .B2(n172), .ZN(
        n127) );
  INV_X1 U207 ( .A(n126), .ZN(n215) );
  AOI22_X1 U208 ( .A1(MVP0[6]), .A2(n142), .B1(eMV0_in[6]), .B2(n172), .ZN(
        n126) );
  INV_X1 U209 ( .A(n125), .ZN(n214) );
  AOI22_X1 U210 ( .A1(MVP0[7]), .A2(n142), .B1(eMV0_in[7]), .B2(n171), .ZN(
        n125) );
  INV_X1 U211 ( .A(n124), .ZN(n213) );
  AOI22_X1 U212 ( .A1(MVP0[8]), .A2(n142), .B1(eMV0_in[8]), .B2(n171), .ZN(
        n124) );
  INV_X1 U213 ( .A(n123), .ZN(n212) );
  AOI22_X1 U214 ( .A1(MVP0[9]), .A2(n142), .B1(eMV0_in[9]), .B2(n170), .ZN(
        n123) );
  INV_X1 U215 ( .A(n132), .ZN(n211) );
  AOI22_X1 U216 ( .A1(MVP0[10]), .A2(n142), .B1(eMV0_in[10]), .B2(n175), .ZN(
        n132) );
  INV_X1 U217 ( .A(n97), .ZN(n197) );
  AOI22_X1 U218 ( .A1(MVP1[13]), .A2(n145), .B1(eMV1_in[13]), .B2(n157), .ZN(
        n97) );
  INV_X1 U219 ( .A(n96), .ZN(n196) );
  AOI22_X1 U220 ( .A1(MVP1[14]), .A2(n145), .B1(eMV1_in[14]), .B2(n157), .ZN(
        n96) );
  INV_X1 U221 ( .A(n95), .ZN(n195) );
  AOI22_X1 U222 ( .A1(MVP1[15]), .A2(n145), .B1(eMV1_in[15]), .B2(n156), .ZN(
        n95) );
  INV_X1 U223 ( .A(n94), .ZN(n194) );
  AOI22_X1 U224 ( .A1(MVP1[16]), .A2(n145), .B1(eMV1_in[16]), .B2(n156), .ZN(
        n94) );
  INV_X1 U225 ( .A(n93), .ZN(n193) );
  AOI22_X1 U226 ( .A1(MVP1[17]), .A2(n145), .B1(eMV1_in[17]), .B2(n155), .ZN(
        n93) );
  INV_X1 U227 ( .A(n92), .ZN(n192) );
  AOI22_X1 U228 ( .A1(MVP1[18]), .A2(n145), .B1(eMV1_in[18]), .B2(n155), .ZN(
        n92) );
  INV_X1 U229 ( .A(n91), .ZN(n191) );
  AOI22_X1 U230 ( .A1(MVP1[19]), .A2(n145), .B1(eMV1_in[19]), .B2(n156), .ZN(
        n91) );
  INV_X1 U231 ( .A(n90), .ZN(n190) );
  AOI22_X1 U232 ( .A1(MVP1[20]), .A2(n145), .B1(eMV1_in[20]), .B2(n155), .ZN(
        n90) );
  INV_X1 U233 ( .A(n78), .ZN(n210) );
  AOI22_X1 U234 ( .A1(MVP2[11]), .A2(n146), .B1(eMV2_in[11]), .B2(n154), .ZN(
        n78) );
  INV_X1 U235 ( .A(n76), .ZN(n209) );
  AOI22_X1 U236 ( .A1(MVP2[12]), .A2(n146), .B1(eMV2_in[12]), .B2(n152), .ZN(
        n76) );
  INV_X1 U237 ( .A(n75), .ZN(n208) );
  AOI22_X1 U238 ( .A1(MVP2[13]), .A2(n146), .B1(eMV2_in[13]), .B2(n151), .ZN(
        n75) );
  INV_X1 U239 ( .A(n74), .ZN(n207) );
  AOI22_X1 U240 ( .A1(MVP2[14]), .A2(n146), .B1(eMV2_in[14]), .B2(n151), .ZN(
        n74) );
  INV_X1 U241 ( .A(n77), .ZN(n200) );
  AOI22_X1 U242 ( .A1(MVP2[21]), .A2(n146), .B1(eMV2_in[21]), .B2(n152), .ZN(
        n77) );
  INV_X1 U243 ( .A(n73), .ZN(n206) );
  AOI22_X1 U244 ( .A1(MVP2[15]), .A2(n147), .B1(eMV2_in[15]), .B2(n150), .ZN(
        n73) );
  INV_X1 U245 ( .A(n72), .ZN(n205) );
  AOI22_X1 U246 ( .A1(MVP2[16]), .A2(n147), .B1(eMV2_in[16]), .B2(n150), .ZN(
        n72) );
  INV_X1 U247 ( .A(n71), .ZN(n204) );
  AOI22_X1 U248 ( .A1(MVP2[17]), .A2(n147), .B1(eMV2_in[17]), .B2(n149), .ZN(
        n71) );
  INV_X1 U249 ( .A(n70), .ZN(n203) );
  AOI22_X1 U250 ( .A1(MVP2[18]), .A2(n147), .B1(eMV2_in[18]), .B2(n149), .ZN(
        n70) );
  INV_X1 U251 ( .A(n69), .ZN(n202) );
  AOI22_X1 U252 ( .A1(MVP2[19]), .A2(n147), .B1(eMV2_in[19]), .B2(n148), .ZN(
        n69) );
  INV_X1 U253 ( .A(n68), .ZN(n201) );
  AOI22_X1 U254 ( .A1(n147), .A2(MVP2[20]), .B1(eMV2_in[20]), .B2(n148), .ZN(
        n68) );
  INV_X1 U255 ( .A(n89), .ZN(n243) );
  AOI22_X1 U256 ( .A1(MVP2[0]), .A2(n145), .B1(eMV2_in[0]), .B2(n154), .ZN(n89) );
  INV_X1 U257 ( .A(n87), .ZN(n242) );
  AOI22_X1 U258 ( .A1(MVP2[1]), .A2(n145), .B1(eMV2_in[1]), .B2(n154), .ZN(n87) );
  INV_X1 U259 ( .A(n86), .ZN(n241) );
  AOI22_X1 U260 ( .A1(MVP2[2]), .A2(n145), .B1(eMV2_in[2]), .B2(n154), .ZN(n86) );
  INV_X1 U261 ( .A(n85), .ZN(n240) );
  AOI22_X1 U262 ( .A1(MVP2[3]), .A2(n146), .B1(eMV2_in[3]), .B2(n153), .ZN(n85) );
  INV_X1 U263 ( .A(n84), .ZN(n239) );
  AOI22_X1 U264 ( .A1(MVP2[4]), .A2(n146), .B1(eMV2_in[4]), .B2(n153), .ZN(n84) );
  INV_X1 U265 ( .A(n83), .ZN(n238) );
  AOI22_X1 U266 ( .A1(MVP2[5]), .A2(n146), .B1(eMV2_in[5]), .B2(n156), .ZN(n83) );
  INV_X1 U267 ( .A(n82), .ZN(n237) );
  AOI22_X1 U268 ( .A1(MVP2[6]), .A2(n146), .B1(eMV2_in[6]), .B2(n155), .ZN(n82) );
  INV_X1 U269 ( .A(n81), .ZN(n236) );
  AOI22_X1 U270 ( .A1(MVP2[7]), .A2(n146), .B1(eMV2_in[7]), .B2(n148), .ZN(n81) );
  INV_X1 U271 ( .A(n80), .ZN(n235) );
  AOI22_X1 U272 ( .A1(MVP2[8]), .A2(n146), .B1(eMV2_in[8]), .B2(n150), .ZN(n80) );
  INV_X1 U273 ( .A(n79), .ZN(n234) );
  AOI22_X1 U274 ( .A1(MVP2[9]), .A2(n146), .B1(eMV2_in[9]), .B2(n153), .ZN(n79) );
  INV_X1 U275 ( .A(n88), .ZN(n233) );
  AOI22_X1 U276 ( .A1(MVP2[10]), .A2(n145), .B1(eMV2_in[10]), .B2(n153), .ZN(
        n88) );
  BUF_X1 U277 ( .A(eIN_SEL), .Z(n140) );
  BUF_X1 U278 ( .A(eIN_SEL), .Z(n141) );
  INV_X1 U280 ( .A(n177), .ZN(n147) );
  INV_X1 U281 ( .A(n135), .ZN(n148) );
  INV_X1 U282 ( .A(n135), .ZN(n149) );
  INV_X1 U283 ( .A(n135), .ZN(n150) );
  INV_X1 U284 ( .A(n135), .ZN(n151) );
  INV_X1 U285 ( .A(n135), .ZN(n152) );
  INV_X1 U286 ( .A(n136), .ZN(n153) );
  INV_X1 U287 ( .A(n136), .ZN(n154) );
  INV_X1 U288 ( .A(n136), .ZN(n155) );
  INV_X1 U289 ( .A(n136), .ZN(n156) );
  INV_X1 U290 ( .A(n137), .ZN(n157) );
  INV_X1 U291 ( .A(n137), .ZN(n158) );
  INV_X1 U292 ( .A(n137), .ZN(n159) );
  INV_X1 U293 ( .A(n137), .ZN(n160) );
  INV_X1 U294 ( .A(n137), .ZN(n161) );
  INV_X1 U295 ( .A(n137), .ZN(n162) );
  INV_X1 U296 ( .A(n137), .ZN(n163) );
  INV_X1 U297 ( .A(n138), .ZN(n164) );
  INV_X1 U298 ( .A(n138), .ZN(n165) );
  INV_X1 U299 ( .A(n138), .ZN(n166) );
  INV_X1 U300 ( .A(n138), .ZN(n167) );
  INV_X1 U301 ( .A(n138), .ZN(n168) );
  INV_X1 U302 ( .A(n138), .ZN(n169) );
  INV_X1 U303 ( .A(n138), .ZN(n170) );
  INV_X1 U304 ( .A(n139), .ZN(n171) );
  INV_X1 U305 ( .A(n139), .ZN(n172) );
  INV_X1 U306 ( .A(n139), .ZN(n173) );
  INV_X1 U307 ( .A(n139), .ZN(n174) );
  INV_X1 U308 ( .A(n139), .ZN(n175) );
  INV_X1 U309 ( .A(n139), .ZN(n176) );
  INV_X1 U310 ( .A(n139), .ZN(n177) );
  INV_X1 constructing_unit_Control_Unit_U22 ( .A(RST), .ZN(
        constructing_unit_Control_Unit_n1) );
  INV_X1 constructing_unit_Control_Unit_U21 ( .A(
        constructing_unit_cmd_SH_EN_int), .ZN(
        constructing_unit_Control_Unit_n6) );
  NOR3_X1 constructing_unit_Control_Unit_U20 ( .A1(
        constructing_unit_Control_Unit_n2), .A2(
        constructing_unit_Control_Unit_n9), .A3(
        constructing_unit_Control_Unit_n8), .ZN(
        constructing_unit_Control_Unit_n11) );
  OAI22_X1 constructing_unit_Control_Unit_U19 ( .A1(
        constructing_unit_Control_Unit_n9), .A2(
        constructing_unit_Control_Unit_n6), .B1(
        constructing_unit_Control_Unit_n11), .B2(
        constructing_unit_Control_Unit_n7), .ZN(
        constructing_unit_Control_Unit_NS[2]) );
  INV_X1 constructing_unit_Control_Unit_U18 ( .A(
        constructing_unit_Control_Unit_START_int), .ZN(
        constructing_unit_Control_Unit_n3) );
  INV_X1 constructing_unit_Control_Unit_U17 ( .A(
        constructing_unit_Control_Unit_GOT_int), .ZN(
        constructing_unit_Control_Unit_n2) );
  AOI22_X1 constructing_unit_Control_Unit_U16 ( .A1(constructing_unit_RST_int), 
        .A2(constructing_unit_Control_Unit_n3), .B1(
        constructing_unit_Control_Unit_PS_1_), .B2(
        constructing_unit_Control_Unit_PS_2_), .ZN(
        constructing_unit_Control_Unit_n16) );
  OAI21_X1 constructing_unit_Control_Unit_U15 ( .B1(
        constructing_unit_Control_Unit_CNT_compEN_OUT_int), .B2(
        constructing_unit_Control_Unit_n7), .A(
        constructing_unit_Control_Unit_n9), .ZN(
        constructing_unit_Control_Unit_n15) );
  OAI211_X1 constructing_unit_Control_Unit_U14 ( .C1(
        constructing_unit_Control_Unit_CNT_STOPcompEN_OUT_int), .C2(
        constructing_unit_Control_Unit_n4), .A(
        constructing_unit_Control_Unit_n15), .B(
        constructing_unit_Control_Unit_n16), .ZN(
        constructing_unit_Control_Unit_NS[0]) );
  NAND2_X1 constructing_unit_Control_Unit_U13 ( .A1(constructing_unit_RST_int), 
        .A2(constructing_unit_Control_Unit_PS_0_), .ZN(
        constructing_unit_Control_Unit_n10) );
  NOR2_X1 constructing_unit_Control_Unit_U12 ( .A1(
        constructing_unit_Control_Unit_n8), .A2(
        constructing_unit_Control_Unit_PS_2_), .ZN(
        constructing_unit_cmd_SH_EN_int) );
  AOI21_X1 constructing_unit_Control_Unit_U11 ( .B1(
        constructing_unit_Control_Unit_PS_2_), .B2(
        constructing_unit_Control_Unit_n2), .A(
        constructing_unit_Control_Unit_n9), .ZN(
        constructing_unit_Control_Unit_n12) );
  OAI221_X1 constructing_unit_Control_Unit_U10 ( .B1(
        constructing_unit_Control_Unit_n12), .B2(
        constructing_unit_Control_Unit_n8), .C1(
        constructing_unit_Control_Unit_n10), .C2(
        constructing_unit_Control_Unit_n3), .A(
        constructing_unit_Control_Unit_n13), .ZN(
        constructing_unit_Control_Unit_NS[1]) );
  NOR2_X1 constructing_unit_Control_Unit_U9 ( .A1(
        constructing_unit_Control_Unit_PS_1_), .A2(
        constructing_unit_Control_Unit_n4), .ZN(cComp_EN) );
  NOR3_X1 constructing_unit_Control_Unit_U8 ( .A1(
        constructing_unit_Control_Unit_n7), .A2(
        constructing_unit_Control_Unit_PS_1_), .A3(
        constructing_unit_Control_Unit_PS_0_), .ZN(
        constructing_unit_CE_compEN_int) );
  NOR2_X1 constructing_unit_Control_Unit_U7 ( .A1(
        constructing_unit_Control_Unit_PS_1_), .A2(
        constructing_unit_Control_Unit_PS_2_), .ZN(constructing_unit_RST_int)
         );
  NOR2_X1 constructing_unit_Control_Unit_U6 ( .A1(
        constructing_unit_Control_Unit_n7), .A2(
        constructing_unit_Control_Unit_n9), .ZN(
        constructing_unit_Control_Unit_n14) );
  NOR2_X1 constructing_unit_Control_Unit_U5 ( .A1(
        constructing_unit_Control_Unit_n4), .A2(
        constructing_unit_Control_Unit_n8), .ZN(cDONE) );
  INV_X1 constructing_unit_Control_Unit_U4 ( .A(
        constructing_unit_Control_Unit_n10), .ZN(cREADY) );
  INV_X1 constructing_unit_Control_Unit_U3 ( .A(
        constructing_unit_Control_Unit_n14), .ZN(
        constructing_unit_Control_Unit_n4) );
  DFFR_X1 constructing_unit_Control_Unit_PS_reg_1_ ( .D(
        constructing_unit_Control_Unit_NS[1]), .CK(clk), .RN(
        constructing_unit_Control_Unit_n1), .Q(
        constructing_unit_Control_Unit_PS_1_), .QN(
        constructing_unit_Control_Unit_n8) );
  DFFR_X1 constructing_unit_Control_Unit_PS_reg_0_ ( .D(
        constructing_unit_Control_Unit_NS[0]), .CK(clk), .RN(
        constructing_unit_Control_Unit_n1), .Q(
        constructing_unit_Control_Unit_PS_0_), .QN(
        constructing_unit_Control_Unit_n9) );
  DFFR_X1 constructing_unit_Control_Unit_PS_reg_2_ ( .D(
        constructing_unit_Control_Unit_NS[2]), .CK(clk), .RN(
        constructing_unit_Control_Unit_n1), .Q(
        constructing_unit_Control_Unit_PS_2_), .QN(
        constructing_unit_Control_Unit_n7) );
  NAND3_X1 constructing_unit_Control_Unit_U23 ( .A1(
        constructing_unit_Control_Unit_n14), .A2(
        constructing_unit_Control_Unit_n8), .A3(
        constructing_unit_Control_Unit_CNT_STOPcompEN_OUT_int), .ZN(
        constructing_unit_Control_Unit_n13) );
  INV_X1 constructing_unit_Control_Unit_START_sampling_U3 ( .A(RST), .ZN(
        constructing_unit_Control_Unit_START_sampling_n1) );
  DFFR_X1 constructing_unit_Control_Unit_START_sampling_Q_int_reg ( .D(START), 
        .CK(clk), .RN(constructing_unit_Control_Unit_START_sampling_n1), .Q(
        constructing_unit_Control_Unit_START_int) );
  INV_X1 constructing_unit_Control_Unit_GOT_sampling_U3 ( .A(RST), .ZN(
        constructing_unit_Control_Unit_GOT_sampling_n1) );
  DFFR_X1 constructing_unit_Control_Unit_GOT_sampling_Q_int_reg ( .D(
        Second_ready), .CK(clk), .RN(
        constructing_unit_Control_Unit_GOT_sampling_n1), .Q(
        constructing_unit_Control_Unit_GOT_int) );
  INV_X1 constructing_unit_Control_Unit_CNT_compEN_OUT_sampling_U3 ( .A(RST), 
        .ZN(constructing_unit_Control_Unit_CNT_compEN_OUT_sampling_n1) );
  DFFR_X1 constructing_unit_Control_Unit_CNT_compEN_OUT_sampling_Q_int_reg ( 
        .D(constructing_unit_CNT_compEN_OUT_int), .CK(clk), .RN(
        constructing_unit_Control_Unit_CNT_compEN_OUT_sampling_n1), .Q(
        constructing_unit_Control_Unit_CNT_compEN_OUT_int) );
  INV_X1 constructing_unit_Control_Unit_CNT_STOPcompEN_OUT_sampling_U3 ( .A(
        RST), .ZN(
        constructing_unit_Control_Unit_CNT_STOPcompEN_OUT_sampling_n1) );
  DFFR_X1 constructing_unit_Control_Unit_CNT_STOPcompEN_OUT_sampling_Q_int_reg ( 
        .D(constructing_unit_CNT_STOPcompEN_OUT_int), .CK(clk), .RN(
        constructing_unit_Control_Unit_CNT_STOPcompEN_OUT_sampling_n1), .Q(
        constructing_unit_Control_Unit_CNT_STOPcompEN_OUT_int) );
  AOI22_X1 constructing_unit_Datapath_U108 ( .A1(
        constructing_unit_Datapath_comp_out_d), .A2(
        constructing_unit_Datapath_D_D_9_), .B1(
        constructing_unit_Datapath_D_min[9]), .B2(
        constructing_unit_Datapath_n2), .ZN(constructing_unit_Datapath_n30) );
  INV_X1 constructing_unit_Datapath_U107 ( .A(constructing_unit_Datapath_n30), 
        .ZN(constructing_unit_Datapath_n67) );
  AOI22_X1 constructing_unit_Datapath_U106 ( .A1(
        constructing_unit_Datapath_D_D_27_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[27]), .B2(
        constructing_unit_Datapath_n4), .ZN(constructing_unit_Datapath_n38) );
  INV_X1 constructing_unit_Datapath_U105 ( .A(constructing_unit_Datapath_n38), 
        .ZN(constructing_unit_Datapath_n21) );
  AOI22_X1 constructing_unit_Datapath_U104 ( .A1(
        constructing_unit_Datapath_D_D_21_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[21]), .B2(
        constructing_unit_Datapath_n6), .ZN(constructing_unit_Datapath_n44) );
  INV_X1 constructing_unit_Datapath_U103 ( .A(constructing_unit_Datapath_n44), 
        .ZN(constructing_unit_Datapath_n27) );
  AOI22_X1 constructing_unit_Datapath_U102 ( .A1(
        constructing_unit_Datapath_D_D_15_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[15]), .B2(
        constructing_unit_Datapath_n9), .ZN(constructing_unit_Datapath_n51) );
  INV_X1 constructing_unit_Datapath_U101 ( .A(constructing_unit_Datapath_n51), 
        .ZN(constructing_unit_Datapath_n61) );
  AOI22_X1 constructing_unit_Datapath_U100 ( .A1(
        constructing_unit_Datapath_D_D_11_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[11]), .B2(
        constructing_unit_Datapath_n10), .ZN(constructing_unit_Datapath_n55)
         );
  INV_X1 constructing_unit_Datapath_U99 ( .A(constructing_unit_Datapath_n55), 
        .ZN(constructing_unit_Datapath_n65) );
  AOI22_X1 constructing_unit_Datapath_U98 ( .A1(
        constructing_unit_Datapath_D_D_23_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[23]), .B2(
        constructing_unit_Datapath_n6), .ZN(constructing_unit_Datapath_n42) );
  INV_X1 constructing_unit_Datapath_U97 ( .A(constructing_unit_Datapath_n42), 
        .ZN(constructing_unit_Datapath_n25) );
  AOI22_X1 constructing_unit_Datapath_U96 ( .A1(
        constructing_unit_Datapath_D_D_17_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[17]), .B2(
        constructing_unit_Datapath_n8), .ZN(constructing_unit_Datapath_n49) );
  INV_X1 constructing_unit_Datapath_U95 ( .A(constructing_unit_Datapath_n49), 
        .ZN(constructing_unit_Datapath_n59) );
  AOI22_X1 constructing_unit_Datapath_U94 ( .A1(
        constructing_unit_Datapath_D_D_19_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[19]), .B2(
        constructing_unit_Datapath_n7), .ZN(constructing_unit_Datapath_n47) );
  INV_X1 constructing_unit_Datapath_U93 ( .A(constructing_unit_Datapath_n47), 
        .ZN(constructing_unit_Datapath_n29) );
  AOI22_X1 constructing_unit_Datapath_U92 ( .A1(
        constructing_unit_Datapath_D_D_13_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[13]), .B2(
        constructing_unit_Datapath_n9), .ZN(constructing_unit_Datapath_n53) );
  INV_X1 constructing_unit_Datapath_U91 ( .A(constructing_unit_Datapath_n53), 
        .ZN(constructing_unit_Datapath_n63) );
  AOI22_X1 constructing_unit_Datapath_U90 ( .A1(
        constructing_unit_Datapath_D_D_5_), .A2(constructing_unit_Datapath_n1), 
        .B1(constructing_unit_Datapath_D_min[5]), .B2(
        constructing_unit_Datapath_n3), .ZN(constructing_unit_Datapath_n34) );
  INV_X1 constructing_unit_Datapath_U89 ( .A(constructing_unit_Datapath_n34), 
        .ZN(constructing_unit_Datapath_n71) );
  AOI22_X1 constructing_unit_Datapath_U88 ( .A1(
        constructing_unit_Datapath_D_D_7_), .A2(constructing_unit_Datapath_n1), 
        .B1(constructing_unit_Datapath_D_min[7]), .B2(
        constructing_unit_Datapath_n2), .ZN(constructing_unit_Datapath_n32) );
  INV_X1 constructing_unit_Datapath_U87 ( .A(constructing_unit_Datapath_n32), 
        .ZN(constructing_unit_Datapath_n69) );
  AOI22_X1 constructing_unit_Datapath_U86 ( .A1(
        constructing_unit_Datapath_D_D_26_), .A2(constructing_unit_Datapath_n1), .B1(constructing_unit_Datapath_D_min[26]), .B2(constructing_unit_Datapath_n5), .ZN(constructing_unit_Datapath_n39) );
  INV_X1 constructing_unit_Datapath_U85 ( .A(constructing_unit_Datapath_n39), 
        .ZN(constructing_unit_Datapath_n22) );
  AOI22_X1 constructing_unit_Datapath_U84 ( .A1(
        constructing_unit_Datapath_D_D_25_), .A2(constructing_unit_Datapath_n1), .B1(constructing_unit_Datapath_D_min[25]), .B2(constructing_unit_Datapath_n5), .ZN(constructing_unit_Datapath_n40) );
  INV_X1 constructing_unit_Datapath_U83 ( .A(constructing_unit_Datapath_n40), 
        .ZN(constructing_unit_Datapath_n23) );
  AOI22_X1 constructing_unit_Datapath_U82 ( .A1(
        constructing_unit_Datapath_D_D_24_), .A2(constructing_unit_Datapath_n1), .B1(constructing_unit_Datapath_D_min[24]), .B2(constructing_unit_Datapath_n5), .ZN(constructing_unit_Datapath_n41) );
  INV_X1 constructing_unit_Datapath_U81 ( .A(constructing_unit_Datapath_n41), 
        .ZN(constructing_unit_Datapath_n24) );
  AOI22_X1 constructing_unit_Datapath_U80 ( .A1(
        constructing_unit_Datapath_D_D_16_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[16]), .B2(
        constructing_unit_Datapath_n8), .ZN(constructing_unit_Datapath_n50) );
  INV_X1 constructing_unit_Datapath_U79 ( .A(constructing_unit_Datapath_n50), 
        .ZN(constructing_unit_Datapath_n60) );
  AOI22_X1 constructing_unit_Datapath_U78 ( .A1(
        constructing_unit_Datapath_D_D_20_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[20]), .B2(
        constructing_unit_Datapath_n7), .ZN(constructing_unit_Datapath_n45) );
  INV_X1 constructing_unit_Datapath_U77 ( .A(constructing_unit_Datapath_n45), 
        .ZN(constructing_unit_Datapath_n28) );
  AOI22_X1 constructing_unit_Datapath_U76 ( .A1(
        constructing_unit_Datapath_D_D_12_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[12]), .B2(
        constructing_unit_Datapath_n10), .ZN(constructing_unit_Datapath_n54)
         );
  INV_X1 constructing_unit_Datapath_U75 ( .A(constructing_unit_Datapath_n54), 
        .ZN(constructing_unit_Datapath_n64) );
  AOI22_X1 constructing_unit_Datapath_U74 ( .A1(
        constructing_unit_Datapath_D_D_22_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[22]), .B2(
        constructing_unit_Datapath_n6), .ZN(constructing_unit_Datapath_n43) );
  INV_X1 constructing_unit_Datapath_U73 ( .A(constructing_unit_Datapath_n43), 
        .ZN(constructing_unit_Datapath_n26) );
  AOI22_X1 constructing_unit_Datapath_U72 ( .A1(
        constructing_unit_Datapath_D_D_18_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[18]), .B2(
        constructing_unit_Datapath_n8), .ZN(constructing_unit_Datapath_n48) );
  INV_X1 constructing_unit_Datapath_U71 ( .A(constructing_unit_Datapath_n48), 
        .ZN(constructing_unit_Datapath_n58) );
  AOI22_X1 constructing_unit_Datapath_U70 ( .A1(
        constructing_unit_Datapath_D_D_14_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[14]), .B2(
        constructing_unit_Datapath_n9), .ZN(constructing_unit_Datapath_n52) );
  INV_X1 constructing_unit_Datapath_U69 ( .A(constructing_unit_Datapath_n52), 
        .ZN(constructing_unit_Datapath_n62) );
  AOI22_X1 constructing_unit_Datapath_U68 ( .A1(
        constructing_unit_Datapath_D_D_10_), .A2(
        constructing_unit_Datapath_comp_out_d), .B1(
        constructing_unit_Datapath_D_min[10]), .B2(
        constructing_unit_Datapath_n10), .ZN(constructing_unit_Datapath_n56)
         );
  INV_X1 constructing_unit_Datapath_U67 ( .A(constructing_unit_Datapath_n56), 
        .ZN(constructing_unit_Datapath_n66) );
  AOI22_X1 constructing_unit_Datapath_U66 ( .A1(
        constructing_unit_Datapath_D_D_2_), .A2(constructing_unit_Datapath_n1), 
        .B1(constructing_unit_Datapath_D_min[2]), .B2(
        constructing_unit_Datapath_n4), .ZN(constructing_unit_Datapath_n37) );
  INV_X1 constructing_unit_Datapath_U65 ( .A(constructing_unit_Datapath_n37), 
        .ZN(constructing_unit_Datapath_n74) );
  AOI22_X1 constructing_unit_Datapath_U64 ( .A1(
        constructing_unit_Datapath_D_D_4_), .A2(constructing_unit_Datapath_n1), 
        .B1(constructing_unit_Datapath_D_min[4]), .B2(
        constructing_unit_Datapath_n3), .ZN(constructing_unit_Datapath_n35) );
  INV_X1 constructing_unit_Datapath_U63 ( .A(constructing_unit_Datapath_n35), 
        .ZN(constructing_unit_Datapath_n72) );
  AOI22_X1 constructing_unit_Datapath_U62 ( .A1(
        constructing_unit_Datapath_D_D_8_), .A2(constructing_unit_Datapath_n1), 
        .B1(constructing_unit_Datapath_D_min[8]), .B2(
        constructing_unit_Datapath_n2), .ZN(constructing_unit_Datapath_n31) );
  INV_X1 constructing_unit_Datapath_U61 ( .A(constructing_unit_Datapath_n31), 
        .ZN(constructing_unit_Datapath_n68) );
  AOI22_X1 constructing_unit_Datapath_U60 ( .A1(
        constructing_unit_Datapath_D_D_6_), .A2(constructing_unit_Datapath_n1), 
        .B1(constructing_unit_Datapath_D_min[6]), .B2(
        constructing_unit_Datapath_n3), .ZN(constructing_unit_Datapath_n33) );
  INV_X1 constructing_unit_Datapath_U59 ( .A(constructing_unit_Datapath_n33), 
        .ZN(constructing_unit_Datapath_n70) );
  BUF_X1 constructing_unit_Datapath_U58 ( .A(
        constructing_unit_Datapath_UA_flag_int_10_), .Z(
        constructing_unit_Datapath_n15) );
  INV_X1 constructing_unit_Datapath_U57 ( .A(
        constructing_unit_Datapath_comp_out_d), .ZN(
        constructing_unit_Datapath_n12) );
  BUF_X1 constructing_unit_Datapath_U56 ( .A(
        constructing_unit_Datapath_UA_flag_int_10_), .Z(
        constructing_unit_Datapath_n14) );
  BUF_X1 constructing_unit_Datapath_U55 ( .A(
        constructing_unit_Datapath_UA_flag_int_10_), .Z(
        constructing_unit_Datapath_n13) );
  AOI22_X1 constructing_unit_Datapath_U54 ( .A1(
        constructing_unit_Datapath_D_D_0_), .A2(constructing_unit_Datapath_n1), 
        .B1(constructing_unit_Datapath_D_min[0]), .B2(
        constructing_unit_Datapath_n11), .ZN(constructing_unit_Datapath_n57)
         );
  AOI22_X1 constructing_unit_Datapath_U53 ( .A1(
        constructing_unit_Datapath_D_D_3_), .A2(constructing_unit_Datapath_n1), 
        .B1(constructing_unit_Datapath_D_min[3]), .B2(
        constructing_unit_Datapath_n4), .ZN(constructing_unit_Datapath_n36) );
  INV_X1 constructing_unit_Datapath_U52 ( .A(constructing_unit_Datapath_n36), 
        .ZN(constructing_unit_Datapath_n73) );
  INV_X1 constructing_unit_Datapath_U51 ( .A(constructing_unit_Datapath_n57), 
        .ZN(constructing_unit_Datapath_n76) );
  AOI22_X1 constructing_unit_Datapath_U50 ( .A1(
        constructing_unit_Datapath_D_D_1_), .A2(constructing_unit_Datapath_n1), 
        .B1(constructing_unit_Datapath_D_min[1]), .B2(
        constructing_unit_Datapath_n7), .ZN(constructing_unit_Datapath_n46) );
  INV_X1 constructing_unit_Datapath_U49 ( .A(constructing_unit_Datapath_n46), 
        .ZN(constructing_unit_Datapath_n75) );
  OR2_X1 constructing_unit_Datapath_U48 ( .A1(
        constructing_unit_Datapath_D_sq[27]), .A2(
        constructing_unit_Datapath_n14), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[27]) );
  BUF_X1 constructing_unit_Datapath_U47 ( .A(
        constructing_unit_Datapath_D_v_14_), .Z(constructing_unit_Datapath_n16) );
  BUF_X1 constructing_unit_Datapath_U46 ( .A(
        constructing_unit_Datapath_D_h_14_), .Z(constructing_unit_Datapath_n17) );
  BUF_X2 constructing_unit_Datapath_U45 ( .A(constructing_unit_RST_int), .Z(
        constructing_unit_Datapath_n20) );
  BUF_X2 constructing_unit_Datapath_U44 ( .A(constructing_unit_RST_int), .Z(
        constructing_unit_Datapath_n19) );
  OR2_X1 constructing_unit_Datapath_U43 ( .A1(
        constructing_unit_Datapath_D_sq[7]), .A2(
        constructing_unit_Datapath_n15), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[7]) );
  OR2_X1 constructing_unit_Datapath_U42 ( .A1(
        constructing_unit_Datapath_D_sq[6]), .A2(
        constructing_unit_Datapath_n15), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[6]) );
  OR2_X1 constructing_unit_Datapath_U41 ( .A1(
        constructing_unit_Datapath_D_sq[5]), .A2(
        constructing_unit_Datapath_n14), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[5]) );
  OR2_X1 constructing_unit_Datapath_U40 ( .A1(
        constructing_unit_Datapath_D_sq[4]), .A2(
        constructing_unit_Datapath_n14), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[4]) );
  OR2_X1 constructing_unit_Datapath_U39 ( .A1(
        constructing_unit_Datapath_D_sq[3]), .A2(
        constructing_unit_Datapath_n14), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[3]) );
  OR2_X1 constructing_unit_Datapath_U38 ( .A1(
        constructing_unit_Datapath_D_sq[2]), .A2(
        constructing_unit_Datapath_n14), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[2]) );
  OR2_X1 constructing_unit_Datapath_U37 ( .A1(
        constructing_unit_Datapath_D_sq[1]), .A2(
        constructing_unit_Datapath_n13), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[1]) );
  OR3_X1 constructing_unit_Datapath_U36 ( .A1(
        constructing_unit_Datapath_UA_flag[2]), .A2(
        constructing_unit_Datapath_UA_flag[1]), .A3(
        constructing_unit_Datapath_UA_flag[0]), .ZN(
        constructing_unit_Datapath_UA_flag_int_0_) );
  BUF_X1 constructing_unit_Datapath_U35 ( .A(constructing_unit_Datapath_n9), 
        .Z(constructing_unit_Datapath_n4) );
  BUF_X1 constructing_unit_Datapath_U34 ( .A(constructing_unit_Datapath_n12), 
        .Z(constructing_unit_Datapath_n5) );
  BUF_X1 constructing_unit_Datapath_U33 ( .A(constructing_unit_Datapath_n2), 
        .Z(constructing_unit_Datapath_n6) );
  BUF_X1 constructing_unit_Datapath_U32 ( .A(constructing_unit_Datapath_n12), 
        .Z(constructing_unit_Datapath_n8) );
  BUF_X1 constructing_unit_Datapath_U31 ( .A(constructing_unit_Datapath_n12), 
        .Z(constructing_unit_Datapath_n10) );
  BUF_X1 constructing_unit_Datapath_U30 ( .A(constructing_unit_Datapath_n12), 
        .Z(constructing_unit_Datapath_n3) );
  BUF_X1 constructing_unit_Datapath_U29 ( .A(constructing_unit_Datapath_n10), 
        .Z(constructing_unit_Datapath_n7) );
  BUF_X1 constructing_unit_Datapath_U28 ( .A(constructing_unit_Datapath_n12), 
        .Z(constructing_unit_Datapath_n9) );
  BUF_X1 constructing_unit_Datapath_U27 ( .A(constructing_unit_Datapath_n12), 
        .Z(constructing_unit_Datapath_n2) );
  OR2_X1 constructing_unit_Datapath_U26 ( .A1(
        constructing_unit_Datapath_D_sq[9]), .A2(
        constructing_unit_Datapath_n15), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[9]) );
  OR2_X1 constructing_unit_Datapath_U25 ( .A1(
        constructing_unit_Datapath_D_sq[8]), .A2(
        constructing_unit_Datapath_n15), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[8]) );
  OR2_X1 constructing_unit_Datapath_U24 ( .A1(
        constructing_unit_Datapath_D_sq[18]), .A2(
        constructing_unit_Datapath_n13), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[18]) );
  OR2_X1 constructing_unit_Datapath_U23 ( .A1(
        constructing_unit_Datapath_D_sq[17]), .A2(
        constructing_unit_Datapath_n13), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[17]) );
  OR2_X1 constructing_unit_Datapath_U22 ( .A1(
        constructing_unit_Datapath_D_sq[16]), .A2(
        constructing_unit_Datapath_n13), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[16]) );
  OR2_X1 constructing_unit_Datapath_U21 ( .A1(
        constructing_unit_Datapath_D_sq[15]), .A2(
        constructing_unit_Datapath_n13), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[15]) );
  OR2_X1 constructing_unit_Datapath_U20 ( .A1(
        constructing_unit_Datapath_D_sq[14]), .A2(
        constructing_unit_Datapath_n13), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[14]) );
  OR2_X1 constructing_unit_Datapath_U19 ( .A1(
        constructing_unit_Datapath_D_sq[13]), .A2(
        constructing_unit_Datapath_n13), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[13]) );
  OR2_X1 constructing_unit_Datapath_U18 ( .A1(
        constructing_unit_Datapath_D_sq[12]), .A2(
        constructing_unit_Datapath_n13), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[12]) );
  OR2_X1 constructing_unit_Datapath_U17 ( .A1(
        constructing_unit_Datapath_D_sq[11]), .A2(
        constructing_unit_Datapath_n13), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[11]) );
  OR2_X1 constructing_unit_Datapath_U16 ( .A1(
        constructing_unit_Datapath_D_sq[10]), .A2(
        constructing_unit_Datapath_n13), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[10]) );
  BUF_X1 constructing_unit_Datapath_U15 ( .A(constructing_unit_Datapath_n12), 
        .Z(constructing_unit_Datapath_n11) );
  AND2_X1 constructing_unit_Datapath_U14 ( .A1(
        constructing_unit_Datapath_comp_out_tmp), .A2(cComp_EN), .ZN(
        constructing_unit_Datapath_comp_out) );
  OR2_X1 constructing_unit_Datapath_U13 ( .A1(
        constructing_unit_Datapath_D_sq[26]), .A2(
        constructing_unit_Datapath_n14), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[26]) );
  OR2_X1 constructing_unit_Datapath_U12 ( .A1(
        constructing_unit_Datapath_D_sq[25]), .A2(
        constructing_unit_Datapath_n14), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[25]) );
  OR2_X1 constructing_unit_Datapath_U11 ( .A1(
        constructing_unit_Datapath_D_sq[24]), .A2(
        constructing_unit_Datapath_n14), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[24]) );
  OR2_X1 constructing_unit_Datapath_U10 ( .A1(
        constructing_unit_Datapath_D_sq[23]), .A2(
        constructing_unit_Datapath_n14), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[23]) );
  OR2_X1 constructing_unit_Datapath_U9 ( .A1(
        constructing_unit_Datapath_D_sq[22]), .A2(
        constructing_unit_Datapath_n14), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[22]) );
  OR2_X1 constructing_unit_Datapath_U8 ( .A1(
        constructing_unit_Datapath_D_sq[21]), .A2(
        constructing_unit_Datapath_n14), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[21]) );
  OR2_X1 constructing_unit_Datapath_U7 ( .A1(
        constructing_unit_Datapath_D_sq[20]), .A2(
        constructing_unit_Datapath_n14), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[20]) );
  OR2_X1 constructing_unit_Datapath_U6 ( .A1(
        constructing_unit_Datapath_D_sq[19]), .A2(
        constructing_unit_Datapath_n13), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[19]) );
  INV_X1 constructing_unit_Datapath_U5 ( .A(constructing_unit_Datapath_n11), 
        .ZN(constructing_unit_Datapath_n1) );
  BUF_X2 constructing_unit_Datapath_U4 ( .A(constructing_unit_RST_int), .Z(
        constructing_unit_Datapath_n18) );
  OR2_X1 constructing_unit_Datapath_U3 ( .A1(
        constructing_unit_Datapath_D_sq[0]), .A2(
        constructing_unit_Datapath_n13), .ZN(
        constructing_unit_Datapath_D_Cur_tmp[0]) );
  INV_X1 constructing_unit_Datapath_L_sub1_sub_19_U14 ( .A(
        constructing_unit_Datapath_MV0_int_v_1__10_), .ZN(
        constructing_unit_Datapath_L_sub1_sub_19_n2) );
  XNOR2_X1 constructing_unit_Datapath_L_sub1_sub_19_U13 ( .A(
        constructing_unit_Datapath_L_sub1_sub_19_n12), .B(
        constructing_unit_Datapath_MV1_int_v_1__0_), .ZN(
        constructing_unit_Datapath_mv1v_mv0v_int[0]) );
  INV_X1 constructing_unit_Datapath_L_sub1_sub_19_U12 ( .A(
        constructing_unit_Datapath_MV0_int_v_1__0_), .ZN(
        constructing_unit_Datapath_L_sub1_sub_19_n12) );
  INV_X1 constructing_unit_Datapath_L_sub1_sub_19_U11 ( .A(
        constructing_unit_Datapath_MV0_int_v_1__9_), .ZN(
        constructing_unit_Datapath_L_sub1_sub_19_n3) );
  INV_X1 constructing_unit_Datapath_L_sub1_sub_19_U10 ( .A(
        constructing_unit_Datapath_MV0_int_v_1__8_), .ZN(
        constructing_unit_Datapath_L_sub1_sub_19_n4) );
  INV_X1 constructing_unit_Datapath_L_sub1_sub_19_U9 ( .A(
        constructing_unit_Datapath_MV0_int_v_1__7_), .ZN(
        constructing_unit_Datapath_L_sub1_sub_19_n5) );
  INV_X1 constructing_unit_Datapath_L_sub1_sub_19_U8 ( .A(
        constructing_unit_Datapath_MV0_int_v_1__6_), .ZN(
        constructing_unit_Datapath_L_sub1_sub_19_n6) );
  INV_X1 constructing_unit_Datapath_L_sub1_sub_19_U7 ( .A(
        constructing_unit_Datapath_MV0_int_v_1__5_), .ZN(
        constructing_unit_Datapath_L_sub1_sub_19_n7) );
  INV_X1 constructing_unit_Datapath_L_sub1_sub_19_U6 ( .A(
        constructing_unit_Datapath_MV0_int_v_1__4_), .ZN(
        constructing_unit_Datapath_L_sub1_sub_19_n8) );
  INV_X1 constructing_unit_Datapath_L_sub1_sub_19_U5 ( .A(
        constructing_unit_Datapath_MV0_int_v_1__3_), .ZN(
        constructing_unit_Datapath_L_sub1_sub_19_n9) );
  INV_X1 constructing_unit_Datapath_L_sub1_sub_19_U4 ( .A(
        constructing_unit_Datapath_MV0_int_v_1__2_), .ZN(
        constructing_unit_Datapath_L_sub1_sub_19_n10) );
  INV_X1 constructing_unit_Datapath_L_sub1_sub_19_U3 ( .A(
        constructing_unit_Datapath_MV1_int_v_1__0_), .ZN(
        constructing_unit_Datapath_L_sub1_sub_19_n1) );
  NAND2_X1 constructing_unit_Datapath_L_sub1_sub_19_U2 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__0_), .A2(
        constructing_unit_Datapath_L_sub1_sub_19_n1), .ZN(
        constructing_unit_Datapath_L_sub1_sub_19_carry[1]) );
  INV_X1 constructing_unit_Datapath_L_sub1_sub_19_U1 ( .A(
        constructing_unit_Datapath_MV0_int_v_1__1_), .ZN(
        constructing_unit_Datapath_L_sub1_sub_19_n11) );
  FA_X1 constructing_unit_Datapath_L_sub1_sub_19_U2_1 ( .A(
        constructing_unit_Datapath_MV1_int_v_1__1_), .B(
        constructing_unit_Datapath_L_sub1_sub_19_n11), .CI(
        constructing_unit_Datapath_L_sub1_sub_19_carry[1]), .CO(
        constructing_unit_Datapath_L_sub1_sub_19_carry[2]), .S(
        constructing_unit_Datapath_mv1v_mv0v_int[1]) );
  FA_X1 constructing_unit_Datapath_L_sub1_sub_19_U2_2 ( .A(
        constructing_unit_Datapath_MV1_int_v_1__2_), .B(
        constructing_unit_Datapath_L_sub1_sub_19_n10), .CI(
        constructing_unit_Datapath_L_sub1_sub_19_carry[2]), .CO(
        constructing_unit_Datapath_L_sub1_sub_19_carry[3]), .S(
        constructing_unit_Datapath_mv1v_mv0v_int[2]) );
  FA_X1 constructing_unit_Datapath_L_sub1_sub_19_U2_3 ( .A(
        constructing_unit_Datapath_MV1_int_v_1__3_), .B(
        constructing_unit_Datapath_L_sub1_sub_19_n9), .CI(
        constructing_unit_Datapath_L_sub1_sub_19_carry[3]), .CO(
        constructing_unit_Datapath_L_sub1_sub_19_carry[4]), .S(
        constructing_unit_Datapath_mv1v_mv0v_int[3]) );
  FA_X1 constructing_unit_Datapath_L_sub1_sub_19_U2_4 ( .A(
        constructing_unit_Datapath_MV1_int_v_1__4_), .B(
        constructing_unit_Datapath_L_sub1_sub_19_n8), .CI(
        constructing_unit_Datapath_L_sub1_sub_19_carry[4]), .CO(
        constructing_unit_Datapath_L_sub1_sub_19_carry[5]), .S(
        constructing_unit_Datapath_mv1v_mv0v_int[4]) );
  FA_X1 constructing_unit_Datapath_L_sub1_sub_19_U2_5 ( .A(
        constructing_unit_Datapath_MV1_int_v_1__5_), .B(
        constructing_unit_Datapath_L_sub1_sub_19_n7), .CI(
        constructing_unit_Datapath_L_sub1_sub_19_carry[5]), .CO(
        constructing_unit_Datapath_L_sub1_sub_19_carry[6]), .S(
        constructing_unit_Datapath_mv1v_mv0v_int[5]) );
  FA_X1 constructing_unit_Datapath_L_sub1_sub_19_U2_6 ( .A(
        constructing_unit_Datapath_MV1_int_v_1__6_), .B(
        constructing_unit_Datapath_L_sub1_sub_19_n6), .CI(
        constructing_unit_Datapath_L_sub1_sub_19_carry[6]), .CO(
        constructing_unit_Datapath_L_sub1_sub_19_carry[7]), .S(
        constructing_unit_Datapath_mv1v_mv0v_int[6]) );
  FA_X1 constructing_unit_Datapath_L_sub1_sub_19_U2_7 ( .A(
        constructing_unit_Datapath_MV1_int_v_1__7_), .B(
        constructing_unit_Datapath_L_sub1_sub_19_n5), .CI(
        constructing_unit_Datapath_L_sub1_sub_19_carry[7]), .CO(
        constructing_unit_Datapath_L_sub1_sub_19_carry[8]), .S(
        constructing_unit_Datapath_mv1v_mv0v_int[7]) );
  FA_X1 constructing_unit_Datapath_L_sub1_sub_19_U2_8 ( .A(
        constructing_unit_Datapath_MV1_int_v_1__8_), .B(
        constructing_unit_Datapath_L_sub1_sub_19_n4), .CI(
        constructing_unit_Datapath_L_sub1_sub_19_carry[8]), .CO(
        constructing_unit_Datapath_L_sub1_sub_19_carry[9]), .S(
        constructing_unit_Datapath_mv1v_mv0v_int[8]) );
  FA_X1 constructing_unit_Datapath_L_sub1_sub_19_U2_9 ( .A(
        constructing_unit_Datapath_MV1_int_v_1__9_), .B(
        constructing_unit_Datapath_L_sub1_sub_19_n3), .CI(
        constructing_unit_Datapath_L_sub1_sub_19_carry[9]), .CO(
        constructing_unit_Datapath_L_sub1_sub_19_carry[10]), .S(
        constructing_unit_Datapath_mv1v_mv0v_int[9]) );
  FA_X1 constructing_unit_Datapath_L_sub1_sub_19_U2_10 ( .A(
        constructing_unit_Datapath_MV1_int_v_1__10_), .B(
        constructing_unit_Datapath_L_sub1_sub_19_n2), .CI(
        constructing_unit_Datapath_L_sub1_sub_19_carry[10]), .CO(
        constructing_unit_Datapath_L_sub1_sub_19_carry[11]), .S(
        constructing_unit_Datapath_mv1v_mv0v_int[10]) );
  FA_X1 constructing_unit_Datapath_L_sub1_sub_19_U2_11 ( .A(
        constructing_unit_Datapath_MV1_int_v_1__10_), .B(
        constructing_unit_Datapath_L_sub1_sub_19_n2), .CI(
        constructing_unit_Datapath_L_sub1_sub_19_carry[11]), .S(
        constructing_unit_Datapath_mv1v_mv0v_int[11]) );
  INV_X1 constructing_unit_Datapath_mv1v_mv0v_REG_0_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_mv1v_mv0v_REG_0_n1) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_0_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[11]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[23]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_0_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[10]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[22]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_0_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[9]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[21]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_0_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[8]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[20]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_0_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[7]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[19]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_0_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[6]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[18]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_0_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[5]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[17]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_0_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[4]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[16]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_0_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[3]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[15]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_0_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[2]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[14]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_0_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[1]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[13]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_0_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[0]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[12]) );
  INV_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_2_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_2_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[12]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[24]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_2_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[13]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[25]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_2_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[14]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[26]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_2_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[15]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[27]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_2_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[16]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[28]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_2_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[17]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[29]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_2_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[18]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[30]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_2_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[19]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[31]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_2_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[20]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[32]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_2_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[21]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[33]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_2_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[22]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[34]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_2_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[23]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[35]) );
  INV_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_3_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_3_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[24]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[36]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_3_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[25]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[37]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_3_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[26]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[38]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_3_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[27]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[39]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_3_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[28]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[40]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_3_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[29]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[41]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_3_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[30]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[42]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_3_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[31]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[43]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_3_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[32]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[44]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_3_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[33]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[45]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_3_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[34]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[46]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_3_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[35]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[47]) );
  INV_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_4_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_4_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[36]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[48]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_4_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[37]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[49]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_4_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[38]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[50]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_4_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[39]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[51]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_4_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[40]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[52]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_4_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[41]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[53]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_4_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[42]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[54]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_4_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[43]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[55]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_4_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[44]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[56]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_4_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[45]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[57]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_4_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[46]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[58]) );
  DFFR_X1 constructing_unit_Datapath_mv1v_mv0v_REG_X_4_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_mv1v_mv0v_int[47]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1v_mv0v_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1v_mv0v_int[59]) );
  INV_X1 constructing_unit_Datapath_h_sample_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_h_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_h_sample_Q_int_reg_0_ ( .D(CU_h[5]), .CK(
        clk), .RN(constructing_unit_Datapath_h_sample_n1), .Q(
        constructing_unit_Datapath_CU_h_int[0]) );
  DFFR_X1 constructing_unit_Datapath_h_sample_Q_int_reg_1_ ( .D(CU_h[6]), .CK(
        clk), .RN(constructing_unit_Datapath_h_sample_n1), .Q(
        constructing_unit_Datapath_CU_h_int[1]) );
  INV_X1 constructing_unit_Datapath_w_sample_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_w_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_w_sample_Q_int_reg_0_ ( .D(CU_w[5]), .CK(
        clk), .RN(constructing_unit_Datapath_w_sample_n1), .Q(
        constructing_unit_Datapath_CU_w_int[0]) );
  DFFR_X1 constructing_unit_Datapath_w_sample_Q_int_reg_1_ ( .D(CU_w[6]), .CK(
        clk), .RN(constructing_unit_Datapath_w_sample_n1), .Q(
        constructing_unit_Datapath_CU_w_int[1]) );
  OR2_X1 constructing_unit_Datapath_hOw_U14 ( .A1(
        constructing_unit_Datapath_hOw_cmd_1_), .A2(
        constructing_unit_Datapath_hOw_n10), .ZN(
        constructing_unit_Datapath_hOw_RSH_in[1]) );
  INV_X1 constructing_unit_Datapath_hOw_U13 ( .A(
        constructing_unit_Datapath_CU_w_int[0]), .ZN(
        constructing_unit_Datapath_hOw_n2) );
  NAND2_X1 constructing_unit_Datapath_hOw_U12 ( .A1(
        constructing_unit_Datapath_CU_w_int[1]), .A2(
        constructing_unit_Datapath_hOw_n3), .ZN(
        constructing_unit_Datapath_hOw_n12) );
  INV_X1 constructing_unit_Datapath_hOw_U11 ( .A(
        constructing_unit_Datapath_CU_h_int[0]), .ZN(
        constructing_unit_Datapath_hOw_n4) );
  INV_X1 constructing_unit_Datapath_hOw_U10 ( .A(
        constructing_unit_Datapath_CU_h_int[1]), .ZN(
        constructing_unit_Datapath_hOw_n3) );
  OR2_X1 constructing_unit_Datapath_hOw_U9 ( .A1(
        constructing_unit_Datapath_hOw_cmd_RSH_out[0]), .A2(
        constructing_unit_Datapath_hOw_cmd_RSH_out[1]), .ZN(
        constructing_unit_Datapath_hOw_RSH_SH_en) );
  OAI21_X1 constructing_unit_Datapath_hOw_U8 ( .B1(
        constructing_unit_Datapath_CU_w_int[1]), .B2(
        constructing_unit_Datapath_hOw_n3), .A(
        constructing_unit_Datapath_hOw_n12), .ZN(
        constructing_unit_Datapath_hOw_n10) );
  NOR2_X1 constructing_unit_Datapath_hOw_U7 ( .A1(
        constructing_unit_Datapath_CU_w_int[0]), .A2(
        constructing_unit_Datapath_hOw_n4), .ZN(
        constructing_unit_Datapath_hOw_n11) );
  OAI21_X1 constructing_unit_Datapath_hOw_U6 ( .B1(
        constructing_unit_Datapath_hOw_n11), .B2(
        constructing_unit_Datapath_hOw_n10), .A(
        constructing_unit_Datapath_hOw_n12), .ZN(
        constructing_unit_Datapath_hOw_n9) );
  INV_X1 constructing_unit_Datapath_hOw_U5 ( .A(
        constructing_unit_Datapath_hOw_n9), .ZN(
        constructing_unit_Datapath_hOw_n1) );
  NOR2_X1 constructing_unit_Datapath_hOw_U4 ( .A1(
        constructing_unit_Datapath_hOw_n3), .A2(
        constructing_unit_Datapath_hOw_n10), .ZN(
        constructing_unit_Datapath_hOw_cmd_1_) );
  OAI22_X1 constructing_unit_Datapath_hOw_U3 ( .A1(
        constructing_unit_Datapath_hOw_n9), .A2(
        constructing_unit_Datapath_hOw_n2), .B1(
        constructing_unit_Datapath_hOw_n1), .B2(
        constructing_unit_Datapath_hOw_n4), .ZN(
        constructing_unit_Datapath_hOw_cmd_0_) );
  OAI22_X1 constructing_unit_Datapath_hOw_U2 ( .A1(
        constructing_unit_Datapath_hOw_n4), .A2(
        constructing_unit_Datapath_hOw_n9), .B1(
        constructing_unit_Datapath_hOw_n1), .B2(
        constructing_unit_Datapath_hOw_n2), .ZN(
        constructing_unit_Datapath_hOw_RSH_in[0]) );
  INV_X1 constructing_unit_Datapath_hOw_FF_X_1_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_hOw_FF_X_1_n1) );
  DFFR_X1 constructing_unit_Datapath_hOw_FF_X_1_Q_int_reg ( .D(
        constructing_unit_Datapath_hOw_n1), .CK(clk), .RN(
        constructing_unit_Datapath_hOw_FF_X_1_n1), .Q(
        constructing_unit_Datapath_hOw_shift_dir_int[1]) );
  INV_X1 constructing_unit_Datapath_hOw_FF_X_2_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_hOw_FF_X_2_n1) );
  DFFR_X1 constructing_unit_Datapath_hOw_FF_X_2_Q_int_reg ( .D(
        constructing_unit_Datapath_hOw_shift_dir_int[1]), .CK(clk), .RN(
        constructing_unit_Datapath_hOw_FF_X_2_n1), .Q(
        constructing_unit_Datapath_hOw_shift_dir_int[2]) );
  INV_X1 constructing_unit_Datapath_hOw_FF_X_3_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_hOw_FF_X_3_n1) );
  DFFR_X1 constructing_unit_Datapath_hOw_FF_X_3_Q_int_reg ( .D(
        constructing_unit_Datapath_hOw_shift_dir_int[2]), .CK(clk), .RN(
        constructing_unit_Datapath_hOw_FF_X_3_n1), .Q(
        constructing_unit_Datapath_SH_cmd_int_2_) );
  INV_X1 constructing_unit_Datapath_hOw_cmd_RSH_U9 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_hOw_cmd_RSH_n2) );
  AOI22_X1 constructing_unit_Datapath_hOw_cmd_RSH_U8 ( .A1(
        constructing_unit_Datapath_hOw_cmd_1_), .A2(cREADY), .B1(
        constructing_unit_Datapath_hOw_cmd_RSH_n4), .B2(
        constructing_unit_Datapath_hOw_cmd_RSH_out[1]), .ZN(
        constructing_unit_Datapath_hOw_cmd_RSH_n7) );
  INV_X1 constructing_unit_Datapath_hOw_cmd_RSH_U7 ( .A(
        constructing_unit_Datapath_hOw_cmd_RSH_n7), .ZN(
        constructing_unit_Datapath_hOw_cmd_RSH_n1) );
  INV_X1 constructing_unit_Datapath_hOw_cmd_RSH_U6 ( .A(cREADY), .ZN(
        constructing_unit_Datapath_hOw_cmd_RSH_n3) );
  AOI22_X1 constructing_unit_Datapath_hOw_cmd_RSH_U5 ( .A1(
        constructing_unit_Datapath_hOw_cmd_RSH_out[1]), .A2(
        constructing_unit_Datapath_hOw_cmd_RSH_n3), .B1(
        constructing_unit_Datapath_hOw_cmd_0_), .B2(cREADY), .ZN(
        constructing_unit_Datapath_hOw_cmd_RSH_n5) );
  NAND2_X1 constructing_unit_Datapath_hOw_cmd_RSH_U4 ( .A1(
        constructing_unit_Datapath_hOw_cmd_RSH_out[0]), .A2(
        constructing_unit_Datapath_hOw_cmd_RSH_n4), .ZN(
        constructing_unit_Datapath_hOw_cmd_RSH_n6) );
  OAI21_X1 constructing_unit_Datapath_hOw_cmd_RSH_U3 ( .B1(
        constructing_unit_Datapath_hOw_cmd_RSH_n4), .B2(
        constructing_unit_Datapath_hOw_cmd_RSH_n5), .A(
        constructing_unit_Datapath_hOw_cmd_RSH_n6), .ZN(
        constructing_unit_Datapath_hOw_cmd_RSH_n8) );
  NOR2_X1 constructing_unit_Datapath_hOw_cmd_RSH_U2 ( .A1(cREADY), .A2(
        constructing_unit_cmd_SH_EN_int), .ZN(
        constructing_unit_Datapath_hOw_cmd_RSH_n4) );
  DFFR_X1 constructing_unit_Datapath_hOw_cmd_RSH_SH_out_int_reg_0_ ( .D(
        constructing_unit_Datapath_hOw_cmd_RSH_n8), .CK(clk), .RN(
        constructing_unit_Datapath_hOw_cmd_RSH_n2), .Q(
        constructing_unit_Datapath_hOw_cmd_RSH_out[0]) );
  DFFR_X1 constructing_unit_Datapath_hOw_cmd_RSH_SH_out_int_reg_1_ ( .D(
        constructing_unit_Datapath_hOw_cmd_RSH_n1), .CK(clk), .RN(
        constructing_unit_Datapath_hOw_cmd_RSH_n2), .Q(
        constructing_unit_Datapath_hOw_cmd_RSH_out[1]) );
  INV_X1 constructing_unit_Datapath_hOw_RSH_U9 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_hOw_RSH_n2) );
  AOI22_X1 constructing_unit_Datapath_hOw_RSH_U8 ( .A1(
        constructing_unit_Datapath_hOw_RSH_in[1]), .A2(cREADY), .B1(
        constructing_unit_Datapath_hOw_RSH_n13), .B2(
        constructing_unit_Datapath_SH_cmd_int_1_), .ZN(
        constructing_unit_Datapath_hOw_RSH_n10) );
  INV_X1 constructing_unit_Datapath_hOw_RSH_U7 ( .A(
        constructing_unit_Datapath_hOw_RSH_n10), .ZN(
        constructing_unit_Datapath_hOw_RSH_n1) );
  INV_X1 constructing_unit_Datapath_hOw_RSH_U6 ( .A(cREADY), .ZN(
        constructing_unit_Datapath_hOw_RSH_n3) );
  AOI22_X1 constructing_unit_Datapath_hOw_RSH_U5 ( .A1(
        constructing_unit_Datapath_SH_cmd_int_1_), .A2(
        constructing_unit_Datapath_hOw_RSH_n3), .B1(
        constructing_unit_Datapath_hOw_RSH_in[0]), .B2(cREADY), .ZN(
        constructing_unit_Datapath_hOw_RSH_n12) );
  NAND2_X1 constructing_unit_Datapath_hOw_RSH_U4 ( .A1(
        constructing_unit_Datapath_SH_cmd_int_0_), .A2(
        constructing_unit_Datapath_hOw_RSH_n13), .ZN(
        constructing_unit_Datapath_hOw_RSH_n11) );
  OAI21_X1 constructing_unit_Datapath_hOw_RSH_U3 ( .B1(
        constructing_unit_Datapath_hOw_RSH_n13), .B2(
        constructing_unit_Datapath_hOw_RSH_n12), .A(
        constructing_unit_Datapath_hOw_RSH_n11), .ZN(
        constructing_unit_Datapath_hOw_RSH_n9) );
  NOR2_X1 constructing_unit_Datapath_hOw_RSH_U2 ( .A1(cREADY), .A2(
        constructing_unit_Datapath_hOw_RSH_SH_en), .ZN(
        constructing_unit_Datapath_hOw_RSH_n13) );
  DFFR_X1 constructing_unit_Datapath_hOw_RSH_SH_out_int_reg_0_ ( .D(
        constructing_unit_Datapath_hOw_RSH_n9), .CK(clk), .RN(
        constructing_unit_Datapath_hOw_RSH_n2), .Q(
        constructing_unit_Datapath_SH_cmd_int_0_) );
  DFFR_X1 constructing_unit_Datapath_hOw_RSH_SH_out_int_reg_1_ ( .D(
        constructing_unit_Datapath_hOw_RSH_n1), .CK(clk), .RN(
        constructing_unit_Datapath_hOw_RSH_n2), .Q(
        constructing_unit_Datapath_SH_cmd_int_1_) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U33 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[13]), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[13]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n26) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U32 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n26), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[13]) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U31 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[12]), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[13]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n27) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U30 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n27), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[12]) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U29 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[11]), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[13]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n28) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U28 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n28), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[11]) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U27 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[10]), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[10]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n29) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U26 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n29), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[10]) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U25 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[8]), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[8]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n18) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U24 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n18), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[8]) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U23 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[7]), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[7]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n19) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U22 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n19), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[7]) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U21 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[6]), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[6]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n20) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U20 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n20), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[6]) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U19 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[5]), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[5]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n21) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U18 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n21), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[5]) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U17 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[4]), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[4]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n22) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U16 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n22), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[4]) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U15 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[3]), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[3]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n23) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U14 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n23), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[3]) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U13 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[2]), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[2]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n24) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U12 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n24), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[2]) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U11 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[1]), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[1]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n25) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U10 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n25), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[1]) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U9 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[0]), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[0]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n30) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U8 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n30), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[0]) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_U7 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .A2(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[9]), .B1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[9]), .B2(
        constructing_unit_Datapath_L_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n17) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U6 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n17), .ZN(
        constructing_unit_Datapath_diff_mult_v_int[9]) );
  OR2_X1 constructing_unit_Datapath_L_LR_SH2_U5 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_shift_amt_int_0_), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_amt_int_1_), .ZN(
        constructing_unit_Datapath_L_LR_SH2_SH_en) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U4 ( .A(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_1_), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n15) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_U3 ( .A(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_), .ZN(
        constructing_unit_Datapath_L_LR_SH2_n16) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_FF_X_1_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_L_LR_SH2_FF_X_1_n1) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_FF_X_1_Q_int_reg ( .D(
        constructing_unit_Datapath_SH_cmd_int_2_), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_FF_X_1_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_1_) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_FF_X_2_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_L_LR_SH2_FF_X_2_n1) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_FF_X_2_Q_int_reg ( .D(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_1_), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_FF_X_2_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_2_) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_FF_X_3_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_L_LR_SH2_FF_X_3_n1) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_FF_X_3_Q_int_reg ( .D(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_2_), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_FF_X_3_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_3_) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_shift_amt_sample_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_L_LR_SH2_shift_amt_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_shift_amt_sample_Q_int_reg_0_ ( 
        .D(constructing_unit_Datapath_SH_cmd_int_0_), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_shift_amt_sample_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_shift_amt_int_0_) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_shift_amt_sample_Q_int_reg_1_ ( 
        .D(constructing_unit_Datapath_SH_cmd_int_1_), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_shift_amt_sample_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_shift_amt_int_1_) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_SH_en2_sampling_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_L_LR_SH2_SH_en2_sampling_n1) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_SH_en2_sampling_Q_int_reg ( .D(
        constructing_unit_Datapath_L_LR_SH2_shift_amt_int_1_), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_SH_en2_sampling_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_SH_en2) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U40 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n1) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U39 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_n15), .A2(
        constructing_unit_Datapath_mv1v_mv0v_int[59]), .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n16), .B2(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[11]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n29) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U38 ( .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n29), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n4) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U37 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[58]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n5) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U36 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[57]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n6) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U35 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[56]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n7) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U34 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[55]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n8) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U33 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[54]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n9) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U32 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[53]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n10) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U31 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[52]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n11) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U30 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[51]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n12) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U29 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[50]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n13) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U28 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[49]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n14) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U27 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[10]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n28) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U26 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[59]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n2) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U25 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n17), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n5), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n18), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n2), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n28), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n40) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U24 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[9]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n27) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U23 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n17), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n6), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n18), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n5), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n27), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n39) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U22 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[8]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n26) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U21 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n17), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n7), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n18), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n6), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n26), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n38) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U20 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[7]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n25) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U19 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n17), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n8), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n18), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n7), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n25), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n37) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U18 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[6]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n24) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U17 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n17), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n9), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n18), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n8), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n24), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n36) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U16 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[5]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n23) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U15 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n17), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n10), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n18), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n9), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n23), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n35) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U14 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[4]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n22) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U13 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n17), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n11), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n18), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n10), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n22), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n34) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U12 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[3]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n21) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U11 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n17), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n12), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n18), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n11), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n21), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n33) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U10 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[2]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n20) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U9 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n17), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n13), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n18), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n12), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n20), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n32) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U8 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[1]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n19) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U7 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n17), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n14), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n18), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n13), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n19), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n31) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U6 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[48]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n15) );
  OAI222_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U5 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n3), .A2(
        constructing_unit_Datapath_L_LR_SH2_n15), .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n15), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n17), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n14), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n18), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n30) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U4 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_SH_en), .A2(
        constructing_unit_Datapath_L_LR_SH2_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n18) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U3 ( .A(
        constructing_unit_Datapath_L_LR_SH2_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n16) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_U2 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_n15), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n18), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n17) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_SH_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_first_n31), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[1]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_SH_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_first_n32), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[2]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_SH_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_first_n33), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[3]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_SH_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_first_n34), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[4]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_SH_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_first_n35), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[5]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_SH_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_first_n36), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[6]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_SH_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_first_n37), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[7]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_SH_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_first_n38), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[8]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_SH_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_first_n39), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[9]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_SH_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_first_n40), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[10]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_SH_out_int_reg_11_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_first_n4), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[11]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_first_SH_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_first_n30), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[0]), .QN(
        constructing_unit_Datapath_L_LR_SH2_RSH_first_n3) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U40 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n1) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U39 ( .A(1'b1), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n16) );
  AOI22_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U38 ( .A1(1'b1), 
        .A2(constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[11]), .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n16), .B2(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[13]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n52) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U37 ( .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n52), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n2) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U36 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[10]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n5) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U35 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[9]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n6) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U34 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[8]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n7) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U33 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[7]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n8) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U32 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[6]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n9) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U31 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[5]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n10) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U30 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[4]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n11) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U29 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[3]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n12) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U28 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[2]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n13) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U27 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[1]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n14) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U26 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[11]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n4) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U25 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[10]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n53) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U24 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n5), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n4), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n53), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n41) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U23 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[9]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n54) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U22 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n6), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n5), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n54), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n42) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U21 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[8]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n55) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U20 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n7), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n6), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n55), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n43) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U19 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[7]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n56) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U18 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n8), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n7), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n56), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n44) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U17 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[6]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n57) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U16 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n9), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n8), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n57), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n45) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U15 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[5]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n58) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U14 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n10), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n9), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n58), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n46) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U13 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[4]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n59) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U12 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n11), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n10), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n59), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n47) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U11 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[3]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n60) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U10 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n12), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n11), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n60), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n48) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U9 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[2]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n61) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U8 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n13), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n12), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n61), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n49) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U7 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[1]), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n62) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U6 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n14), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n13), .A(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n62), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n50) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U5 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1R[0]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n15) );
  OAI222_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U4 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n65), .A2(1'b1), .B1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n15), .B2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n64), .C1(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n14), .C2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n63), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n51) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U3 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_SH_en2), .A2(1'b1), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n63) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_U2 ( .A1(1'b1), .A2(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n63), .ZN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n64) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_SH_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_second_n51), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[0]), .QN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n65) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_SH_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_second_n50), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[1]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_SH_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_second_n49), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[2]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_SH_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_second_n48), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[3]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_SH_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_second_n47), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[4]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_SH_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_second_n46), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[5]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_SH_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_second_n45), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[6]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_SH_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_second_n44), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[7]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_SH_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_second_n43), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[8]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_SH_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_second_n42), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[9]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_SH_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_second_n41), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[10]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_RSH_second_SH_out_int_reg_11_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_RSH_second_n2), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2R_ext[13]) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U42 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U41 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[58]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n4) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U40 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[57]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n5) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U39 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[56]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n6) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U38 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[55]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n7) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U37 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[54]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n8) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U36 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[53]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n9) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U35 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[52]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n10) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U34 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[51]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n11) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U33 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[50]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n12) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U32 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[49]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n13) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U31 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[48]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n14) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U30 ( .A(
        constructing_unit_Datapath_mv1v_mv0v_int[59]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n3) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U29 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[0]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n17) );
  OAI21_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U28 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n16), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n14), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n17), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n30) );
  OAI22_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U27 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n3), .B1(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_1_), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n2), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n42) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U26 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[1]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n19) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U25 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n14), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n18), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n16), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n13), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n19), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n31) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U24 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[11]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n29) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U23 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n18), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n4), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n16), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n3), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n29), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n41) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U22 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[10]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n28) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U21 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n18), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n5), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n16), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n4), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n28), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n40) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U20 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[9]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n27) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U19 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n18), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n6), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n16), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n5), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n27), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n39) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U18 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[8]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n26) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U17 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n18), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n7), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n16), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n6), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n26), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n38) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U16 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[7]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n25) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U15 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n18), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n8), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n16), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n7), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n25), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n37) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U14 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[6]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n24) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U13 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n18), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n9), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n16), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n8), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n24), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n36) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U12 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[5]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n23) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U11 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n18), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n10), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n16), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n9), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n23), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n35) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U10 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[4]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n22) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U9 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n18), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n11), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n16), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n10), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n22), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n34) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U8 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[3]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n21) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U7 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n18), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n12), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n16), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n11), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n21), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n33) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U6 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[2]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n20) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U5 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n18), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n13), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n16), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n12), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n20), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n32) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U4 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_1_), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n18), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n16) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U3 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_SH_en), .A2(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_1_), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n18) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_U2 ( .A(
        constructing_unit_Datapath_L_LR_SH2_shift_dir_int_1_), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n15) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_SH_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_first_n32), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[2]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_SH_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_first_n33), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[3]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_SH_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_first_n34), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[4]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_SH_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_first_n35), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[5]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_SH_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_first_n36), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[6]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_SH_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_first_n37), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[7]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_SH_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_first_n38), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[8]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_SH_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_first_n39), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[9]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_SH_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_first_n40), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[10]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_SH_out_int_reg_11_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_first_n41), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[11]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_SH_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_first_n31), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[1]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_SH_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_first_n30), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[0]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_first_SH_out_int_reg_12_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_first_n42), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[12]), .QN(
        constructing_unit_Datapath_L_LR_SH2_LSH_first_n2) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U45 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U44 ( .A(1'b1), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U43 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[12]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n3) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U42 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[11]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n4) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U41 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[10]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n5) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U40 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[9]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n6) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U39 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[8]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n7) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U38 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[7]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n8) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U37 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[6]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n9) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U36 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[5]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n10) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U35 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[4]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n11) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U34 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[3]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n12) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U33 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[2]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n13) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U32 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[1]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n14) );
  INV_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U31 ( .A(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d1L[0]), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n15) );
  OAI22_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U30 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n3), .B1(1'b1), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n2), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n45) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U29 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[0]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n18) );
  OAI21_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U28 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n15), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n18), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n32) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U27 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[1]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n20) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U26 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n15), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n14), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n20), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n33) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U25 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[12]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n31) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U24 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n4), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n3), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n31), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n44) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U23 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[11]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n30) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U22 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n5), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n4), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n30), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n43) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U21 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[10]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n29) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U20 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n6), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n5), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n29), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n42) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U19 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[9]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n28) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U18 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n7), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n6), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n28), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n41) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U17 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[8]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n27) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U16 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n8), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n7), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n27), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n40) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U15 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[7]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n26) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U14 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n9), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n8), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n26), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n39) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U13 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[6]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n25) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U12 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n10), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n9), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n25), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n38) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U11 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[5]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n24) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U10 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n11), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n10), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n24), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n37) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U9 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[4]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n23) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U8 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n12), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n11), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n23), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n36) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U7 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[3]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n22) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U6 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n13), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n12), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n22), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n35) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U5 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[2]), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n21) );
  OAI221_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U4 ( .B1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19), .B2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n14), .C1(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17), .C2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n13), .A(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n21), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n34) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U3 ( .A1(1'b1), .A2(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n17) );
  NAND2_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_U2 ( .A1(
        constructing_unit_Datapath_L_LR_SH2_SH_en2), .A2(1'b1), .ZN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n19) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n33), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[1]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n34), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[2]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n35), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[3]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n36), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[4]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n37), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[5]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n38), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[6]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n39), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[7]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n40), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[8]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n41), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[9]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n42), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[10]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_11_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n43), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[11]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_12_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n44), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[12]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n32), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[0]) );
  DFFR_X1 constructing_unit_Datapath_L_LR_SH2_LSH_second_SH_out_int_reg_13_ ( 
        .D(constructing_unit_Datapath_L_LR_SH2_LSH_second_n45), .CK(clk), .RN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_L_LR_SH2_MV1_MV0_d2L[13]), .QN(
        constructing_unit_Datapath_L_LR_SH2_LSH_second_n2) );
  INV_X1 constructing_unit_Datapath_diff_mult_v_int_samp_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[0]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[14]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[1]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[15]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[2]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[16]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[3]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[17]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[4]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[18]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[5]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[19]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[6]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[20]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[7]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[21]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[8]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[22]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[10]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[24]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[11]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[25]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[12]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[26]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[13]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[27]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_v_int_samp_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_diff_mult_v_int[9]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_v_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_v_int[23]) );
  INV_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[0]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[11]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[1]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[12]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[2]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[13]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[3]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[14]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[4]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[15]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[5]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[16]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[6]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[17]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[7]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[18]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[8]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[19]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[9]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[20]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[21]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[22]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[23]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_h_ext_sample_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_MV0_int_h_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[24]) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U17 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[27]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n2) );
  XNOR2_X1 constructing_unit_Datapath_L_sub2_sub_19_U16 ( .A(
        constructing_unit_Datapath_L_sub2_sub_19_n15), .B(
        constructing_unit_Datapath_MV0_int_h_ext[11]), .ZN(
        constructing_unit_Datapath_MV2p_int_h[0]) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U15 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[14]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n15) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U14 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[26]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n3) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U13 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[25]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n4) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U12 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[24]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n5) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U11 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[23]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n6) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U10 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[22]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n7) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U9 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[21]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n8) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U8 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[20]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n9) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U7 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[19]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n10) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U6 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[18]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n11) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U5 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[17]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n12) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U4 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[16]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n13) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U3 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[11]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n1) );
  NAND2_X1 constructing_unit_Datapath_L_sub2_sub_19_U2 ( .A1(
        constructing_unit_Datapath_diff_mult_v_int[14]), .A2(
        constructing_unit_Datapath_L_sub2_sub_19_n1), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_carry[1]) );
  INV_X1 constructing_unit_Datapath_L_sub2_sub_19_U1 ( .A(
        constructing_unit_Datapath_diff_mult_v_int[15]), .ZN(
        constructing_unit_Datapath_L_sub2_sub_19_n14) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_1 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[12]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n14), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[1]), .CO(
        constructing_unit_Datapath_L_sub2_sub_19_carry[2]), .S(
        constructing_unit_Datapath_MV2p_int_h[1]) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_2 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[13]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n13), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[2]), .CO(
        constructing_unit_Datapath_L_sub2_sub_19_carry[3]), .S(
        constructing_unit_Datapath_MV2p_int_h[2]) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_3 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[14]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n12), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[3]), .CO(
        constructing_unit_Datapath_L_sub2_sub_19_carry[4]), .S(
        constructing_unit_Datapath_MV2p_int_h[3]) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_4 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[15]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n11), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[4]), .CO(
        constructing_unit_Datapath_L_sub2_sub_19_carry[5]), .S(
        constructing_unit_Datapath_MV2p_int_h[4]) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_5 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[16]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n10), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[5]), .CO(
        constructing_unit_Datapath_L_sub2_sub_19_carry[6]), .S(
        constructing_unit_Datapath_MV2p_int_h[5]) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_6 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[17]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n9), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[6]), .CO(
        constructing_unit_Datapath_L_sub2_sub_19_carry[7]), .S(
        constructing_unit_Datapath_MV2p_int_h[6]) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_7 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[18]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n8), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[7]), .CO(
        constructing_unit_Datapath_L_sub2_sub_19_carry[8]), .S(
        constructing_unit_Datapath_MV2p_int_h[7]) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_8 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[19]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n7), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[8]), .CO(
        constructing_unit_Datapath_L_sub2_sub_19_carry[9]), .S(
        constructing_unit_Datapath_MV2p_int_h[8]) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_9 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[20]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n6), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[9]), .CO(
        constructing_unit_Datapath_L_sub2_sub_19_carry[10]), .S(
        constructing_unit_Datapath_MV2p_int_h[9]) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_10 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[21]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n5), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[10]), .CO(
        constructing_unit_Datapath_L_sub2_sub_19_carry[11]), .S(
        constructing_unit_Datapath_MV2p_int_h[10]) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_11 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[22]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n4), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[11]), .CO(
        constructing_unit_Datapath_L_sub2_sub_19_carry[12]), .S(
        constructing_unit_Datapath_MV2p_int_h[11]) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_12 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[23]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n3), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[12]), .CO(
        constructing_unit_Datapath_L_sub2_sub_19_carry[13]), .S(
        constructing_unit_Datapath_MV2p_int_h[12]) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_13 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[24]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n2), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[13]), .CO(
        constructing_unit_Datapath_L_sub2_sub_19_carry[14]), .S(
        constructing_unit_Datapath_MV2p_int_h[13]) );
  FA_X1 constructing_unit_Datapath_L_sub2_sub_19_U2_14 ( .A(
        constructing_unit_Datapath_MV0_int_h_ext[24]), .B(
        constructing_unit_Datapath_L_sub2_sub_19_n2), .CI(
        constructing_unit_Datapath_L_sub2_sub_19_carry[14]), .S(
        constructing_unit_Datapath_MV2p_int_h[14]) );
  INV_X1 constructing_unit_Datapath_MV2p_int_h_sample_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_14_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[14]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[29]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[13]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[28]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[12]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[27]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[11]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[26]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[25]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[9]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[24]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[8]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[23]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[7]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[22]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[6]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[21]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[5]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[20]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[4]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[19]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[3]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[18]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[2]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[17]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[1]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[16]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_h_sample_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_MV2p_int_h[0]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_h_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_h[15]) );
  INV_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_U4 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n2) );
  INV_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[0]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[11]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[1]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[12]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[2]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[13]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[3]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[14]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[4]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[15]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[5]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[16]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[6]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[17]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[7]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[18]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[8]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[19]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[9]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[20]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[21]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[22]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n2), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[23]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n2), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[24]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_h_ext_sample_Q_int_reg_14_ ( .D(
        constructing_unit_Datapath_MV2_int_h_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_h_ext_sample_n2), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[25]) );
  XNOR2_X1 constructing_unit_Datapath_L_subD_sub_19_U18 ( .A(
        constructing_unit_Datapath_L_subD_sub_19_n16), .B(
        constructing_unit_Datapath_MV2p_int_h[15]), .ZN(
        constructing_unit_Datapath_D_h_tmp[0]) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U17 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[11]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n16) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U16 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[25]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n2) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U15 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[24]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n3) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U14 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[23]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n4) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U13 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[22]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n5) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U12 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[21]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n6) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U11 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[20]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n7) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U10 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[19]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n8) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U9 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[18]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n9) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U8 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[17]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n10) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U7 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[16]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n11) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U6 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[15]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n12) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U5 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[14]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n13) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U4 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[13]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n14) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U3 ( .A(
        constructing_unit_Datapath_MV2p_int_h[15]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n1) );
  NAND2_X1 constructing_unit_Datapath_L_subD_sub_19_U2 ( .A1(
        constructing_unit_Datapath_MV2_int_h_ext[11]), .A2(
        constructing_unit_Datapath_L_subD_sub_19_n1), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_carry[1]) );
  INV_X1 constructing_unit_Datapath_L_subD_sub_19_U1 ( .A(
        constructing_unit_Datapath_MV2_int_h_ext[12]), .ZN(
        constructing_unit_Datapath_L_subD_sub_19_n15) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_1 ( .A(
        constructing_unit_Datapath_MV2p_int_h[16]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n15), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[1]), .CO(
        constructing_unit_Datapath_L_subD_sub_19_carry[2]), .S(
        constructing_unit_Datapath_D_h_tmp[1]) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_2 ( .A(
        constructing_unit_Datapath_MV2p_int_h[17]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n14), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[2]), .CO(
        constructing_unit_Datapath_L_subD_sub_19_carry[3]), .S(
        constructing_unit_Datapath_D_h_tmp[2]) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_3 ( .A(
        constructing_unit_Datapath_MV2p_int_h[18]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n13), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[3]), .CO(
        constructing_unit_Datapath_L_subD_sub_19_carry[4]), .S(
        constructing_unit_Datapath_D_h_tmp[3]) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_4 ( .A(
        constructing_unit_Datapath_MV2p_int_h[19]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n12), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[4]), .CO(
        constructing_unit_Datapath_L_subD_sub_19_carry[5]), .S(
        constructing_unit_Datapath_D_h_tmp[4]) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_5 ( .A(
        constructing_unit_Datapath_MV2p_int_h[20]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n11), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[5]), .CO(
        constructing_unit_Datapath_L_subD_sub_19_carry[6]), .S(
        constructing_unit_Datapath_D_h_tmp[5]) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_6 ( .A(
        constructing_unit_Datapath_MV2p_int_h[21]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n10), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[6]), .CO(
        constructing_unit_Datapath_L_subD_sub_19_carry[7]), .S(
        constructing_unit_Datapath_D_h_tmp[6]) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_7 ( .A(
        constructing_unit_Datapath_MV2p_int_h[22]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n9), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[7]), .CO(
        constructing_unit_Datapath_L_subD_sub_19_carry[8]), .S(
        constructing_unit_Datapath_D_h_tmp[7]) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_8 ( .A(
        constructing_unit_Datapath_MV2p_int_h[23]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n8), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[8]), .CO(
        constructing_unit_Datapath_L_subD_sub_19_carry[9]), .S(
        constructing_unit_Datapath_D_h_tmp[8]) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_9 ( .A(
        constructing_unit_Datapath_MV2p_int_h[24]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n7), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[9]), .CO(
        constructing_unit_Datapath_L_subD_sub_19_carry[10]), .S(
        constructing_unit_Datapath_D_h_tmp[9]) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_10 ( .A(
        constructing_unit_Datapath_MV2p_int_h[25]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n6), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[10]), .CO(
        constructing_unit_Datapath_L_subD_sub_19_carry[11]), .S(
        constructing_unit_Datapath_D_h_tmp[10]) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_11 ( .A(
        constructing_unit_Datapath_MV2p_int_h[26]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n5), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[11]), .CO(
        constructing_unit_Datapath_L_subD_sub_19_carry[12]), .S(
        constructing_unit_Datapath_D_h_tmp[11]) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_12 ( .A(
        constructing_unit_Datapath_MV2p_int_h[27]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n4), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[12]), .CO(
        constructing_unit_Datapath_L_subD_sub_19_carry[13]), .S(
        constructing_unit_Datapath_D_h_tmp[12]) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_13 ( .A(
        constructing_unit_Datapath_MV2p_int_h[28]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n3), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[13]), .CO(
        constructing_unit_Datapath_L_subD_sub_19_carry[14]), .S(
        constructing_unit_Datapath_D_h_tmp[13]) );
  FA_X1 constructing_unit_Datapath_L_subD_sub_19_U2_14 ( .A(
        constructing_unit_Datapath_MV2p_int_h[29]), .B(
        constructing_unit_Datapath_L_subD_sub_19_n2), .CI(
        constructing_unit_Datapath_L_subD_sub_19_carry[14]), .S(
        constructing_unit_Datapath_D_h_tmp[14]) );
  INV_X1 constructing_unit_Datapath_D_h_sample_U4 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_D_h_sample_n2) );
  INV_X1 constructing_unit_Datapath_D_h_sample_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_D_h_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_D_h_tmp[0]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n1), .Q(
        constructing_unit_Datapath_D_h_0_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_D_h_tmp[1]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n1), .Q(
        constructing_unit_Datapath_D_h_1_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_D_h_tmp[2]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n1), .Q(
        constructing_unit_Datapath_D_h_2_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_D_h_tmp[3]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n1), .Q(
        constructing_unit_Datapath_D_h_3_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_D_h_tmp[4]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n1), .Q(
        constructing_unit_Datapath_D_h_4_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_D_h_tmp[5]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n1), .Q(
        constructing_unit_Datapath_D_h_5_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_D_h_tmp[6]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n1), .Q(
        constructing_unit_Datapath_D_h_6_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_D_h_tmp[7]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n1), .Q(
        constructing_unit_Datapath_D_h_7_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_D_h_tmp[8]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n1), .Q(
        constructing_unit_Datapath_D_h_8_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_D_h_tmp[9]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n1), .Q(
        constructing_unit_Datapath_D_h_9_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_D_h_tmp[10]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n1), .Q(
        constructing_unit_Datapath_D_h_10_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_D_h_tmp[11]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n1), .Q(
        constructing_unit_Datapath_D_h_11_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_D_h_tmp[12]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n2), .Q(
        constructing_unit_Datapath_D_h_12_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_D_h_tmp[13]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n2), .Q(
        constructing_unit_Datapath_D_h_13_) );
  DFFR_X1 constructing_unit_Datapath_D_h_sample_Q_int_reg_14_ ( .D(
        constructing_unit_Datapath_D_h_tmp[14]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sample_n2), .Q(
        constructing_unit_Datapath_D_h_14_) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U826 ( .A(
        constructing_unit_Datapath_D_h_13_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n776) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U825 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n666), .B(
        constructing_unit_Datapath_D_h_6_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n848) );
  NAND2_X1 constructing_unit_Datapath_L_squarer_mult_13_U824 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n848), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n763) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U823 ( .A(
        constructing_unit_Datapath_n17), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n778) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U822 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n776), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n778), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n112) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U821 ( .A(
        constructing_unit_Datapath_D_h_13_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n758) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U820 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n664), .B(
        constructing_unit_Datapath_D_h_4_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n847) );
  NAND2_X1 constructing_unit_Datapath_L_squarer_mult_13_U819 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n847), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n745) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U818 ( .A(
        constructing_unit_Datapath_n17), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n760) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U817 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n758), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n760), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n134) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U816 ( .A(
        constructing_unit_Datapath_D_h_13_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n740) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U815 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n662), .B(
        constructing_unit_Datapath_D_h_2_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n846) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U814 ( .A(
        constructing_unit_Datapath_n17), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n742) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U813 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n740), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n742), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n160) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U812 ( .A(
        constructing_unit_Datapath_D_h_2_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n809) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U811 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n672), .B(
        constructing_unit_Datapath_D_h_12_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n845) );
  NAND2_X1 constructing_unit_Datapath_L_squarer_mult_13_U810 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n845), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n706) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U809 ( .A(
        constructing_unit_Datapath_D_h_3_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n810) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U808 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n809), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n810), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n844) );
  XOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U807 ( .A(
        constructing_unit_Datapath_D_h_1_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n674), .Z(
        constructing_unit_Datapath_L_squarer_mult_13_n843) );
  NAND2_X1 constructing_unit_Datapath_L_squarer_mult_13_U806 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n843), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n689), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n842) );
  NAND2_X1 constructing_unit_Datapath_L_squarer_mult_13_U805 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n690), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n842), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n174) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U804 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n842), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n690), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n175) );
  AND3_X1 constructing_unit_Datapath_L_squarer_mult_13_U803 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n674), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n691), .A3(
        constructing_unit_Datapath_L_squarer_mult_13_n689), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n284) );
  OR3_X1 constructing_unit_Datapath_L_squarer_mult_13_U802 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .A2(
        constructing_unit_Datapath_D_h_0_), .A3(
        constructing_unit_Datapath_L_squarer_mult_13_n672), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n841) );
  OAI21_X1 constructing_unit_Datapath_L_squarer_mult_13_U801 ( .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n672), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .A(
        constructing_unit_Datapath_L_squarer_mult_13_n841), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n285) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U800 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n670), .B(
        constructing_unit_Datapath_D_h_10_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n840) );
  NAND2_X1 constructing_unit_Datapath_L_squarer_mult_13_U799 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n840), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n702) );
  OR3_X1 constructing_unit_Datapath_L_squarer_mult_13_U798 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .A2(
        constructing_unit_Datapath_D_h_0_), .A3(
        constructing_unit_Datapath_L_squarer_mult_13_n670), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n839) );
  OAI21_X1 constructing_unit_Datapath_L_squarer_mult_13_U797 ( .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n670), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .A(
        constructing_unit_Datapath_L_squarer_mult_13_n839), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n286) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U796 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n668), .B(
        constructing_unit_Datapath_D_h_8_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n838) );
  NAND2_X1 constructing_unit_Datapath_L_squarer_mult_13_U795 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n838), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n698) );
  OR3_X1 constructing_unit_Datapath_L_squarer_mult_13_U794 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .A2(
        constructing_unit_Datapath_D_h_0_), .A3(
        constructing_unit_Datapath_L_squarer_mult_13_n668), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n837) );
  OAI21_X1 constructing_unit_Datapath_L_squarer_mult_13_U793 ( .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n668), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .A(
        constructing_unit_Datapath_L_squarer_mult_13_n837), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n287) );
  OR3_X1 constructing_unit_Datapath_L_squarer_mult_13_U792 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .A2(
        constructing_unit_Datapath_D_h_0_), .A3(
        constructing_unit_Datapath_L_squarer_mult_13_n666), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n836) );
  OAI21_X1 constructing_unit_Datapath_L_squarer_mult_13_U791 ( .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n666), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .A(
        constructing_unit_Datapath_L_squarer_mult_13_n836), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n288) );
  OR3_X1 constructing_unit_Datapath_L_squarer_mult_13_U790 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .A2(
        constructing_unit_Datapath_D_h_0_), .A3(
        constructing_unit_Datapath_L_squarer_mult_13_n664), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n835) );
  OAI21_X1 constructing_unit_Datapath_L_squarer_mult_13_U789 ( .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n664), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .A(
        constructing_unit_Datapath_L_squarer_mult_13_n835), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n289) );
  OR3_X1 constructing_unit_Datapath_L_squarer_mult_13_U788 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .A2(
        constructing_unit_Datapath_D_h_0_), .A3(
        constructing_unit_Datapath_L_squarer_mult_13_n662), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n834) );
  OAI21_X1 constructing_unit_Datapath_L_squarer_mult_13_U787 ( .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n662), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .A(
        constructing_unit_Datapath_L_squarer_mult_13_n834), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n290) );
  NAND2_X1 constructing_unit_Datapath_L_squarer_mult_13_U786 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n709) );
  OAI21_X1 constructing_unit_Datapath_L_squarer_mult_13_U785 ( .B1(
        constructing_unit_Datapath_D_h_0_), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n660), .A(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n291) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U784 ( .A(
        constructing_unit_Datapath_D_h_13_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n833) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U783 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n833), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n293) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U782 ( .A(
        constructing_unit_Datapath_D_h_12_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n832) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U781 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n832), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n294) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U780 ( .A(
        constructing_unit_Datapath_D_h_11_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n831) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U779 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n831), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n295) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U778 ( .A(
        constructing_unit_Datapath_D_h_10_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n830) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U777 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n830), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n296) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U776 ( .A(
        constructing_unit_Datapath_D_h_9_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n829) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U775 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n829), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n297) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U774 ( .A(
        constructing_unit_Datapath_D_h_8_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n828) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U773 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n828), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n298) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U772 ( .A(
        constructing_unit_Datapath_D_h_7_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n827) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U771 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n827), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n299) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U770 ( .A(
        constructing_unit_Datapath_D_h_6_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n826) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U769 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n826), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n300) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U768 ( .A(
        constructing_unit_Datapath_D_h_5_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n825) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U767 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n825), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n301) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U766 ( .A(
        constructing_unit_Datapath_D_h_4_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n824) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U765 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n824), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n302) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U764 ( .A(
        constructing_unit_Datapath_D_h_3_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n823) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U763 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n823), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n303) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U762 ( .A(
        constructing_unit_Datapath_D_h_2_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n822) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U761 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n822), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n304) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U760 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n691), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n306) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U759 ( .A(
        constructing_unit_Datapath_n17), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n708) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U758 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n708), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n708), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n820) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U757 ( .A(
        constructing_unit_Datapath_D_h_12_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n819) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U756 ( .A(
        constructing_unit_Datapath_D_h_13_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n705) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U755 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n819), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n705), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n308) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U754 ( .A(
        constructing_unit_Datapath_D_h_11_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n818) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U753 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n818), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n819), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n309) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U752 ( .A(
        constructing_unit_Datapath_D_h_10_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n817) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U751 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n817), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n818), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n310) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U750 ( .A(
        constructing_unit_Datapath_D_h_9_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n816) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U749 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n816), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n817), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n311) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U748 ( .A(
        constructing_unit_Datapath_D_h_8_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n815) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U747 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n815), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n816), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n312) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U746 ( .A(
        constructing_unit_Datapath_D_h_7_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n814) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U745 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n814), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n815), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n313) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U744 ( .A(
        constructing_unit_Datapath_D_h_6_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n813) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U743 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n813), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n814), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n314) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U742 ( .A(
        constructing_unit_Datapath_D_h_5_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n812) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U741 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n812), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n813), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n315) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U740 ( .A(
        constructing_unit_Datapath_D_h_4_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n811) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U739 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n811), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n812), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n316) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U738 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n810), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n811), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n317) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U737 ( .A(
        constructing_unit_Datapath_D_h_1_), .B(
        constructing_unit_Datapath_D_h_13_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n808) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U736 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n808), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n809), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n319) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U735 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n671), .B(
        constructing_unit_Datapath_D_h_0_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n807) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U734 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n807), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n808), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n320) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U733 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n691), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n321) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U732 ( .A(
        constructing_unit_Datapath_n17), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n704) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U731 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n704), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n704), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n806) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U730 ( .A(
        constructing_unit_Datapath_D_h_12_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n805) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U729 ( .A(
        constructing_unit_Datapath_D_h_13_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n701) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U728 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n805), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n701), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n323) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U727 ( .A(
        constructing_unit_Datapath_D_h_11_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n804) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U726 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n804), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n805), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n324) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U725 ( .A(
        constructing_unit_Datapath_D_h_10_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n803) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U724 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n803), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n804), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n325) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U723 ( .A(
        constructing_unit_Datapath_D_h_9_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n802) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U722 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n802), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n803), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n326) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U721 ( .A(
        constructing_unit_Datapath_D_h_8_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n801) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U720 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n801), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n802), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n327) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U719 ( .A(
        constructing_unit_Datapath_D_h_7_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n800) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U718 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n800), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n801), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n328) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U717 ( .A(
        constructing_unit_Datapath_D_h_6_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n799) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U716 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n799), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n800), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n329) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U715 ( .A(
        constructing_unit_Datapath_D_h_5_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n798) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U714 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n798), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n799), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n330) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U713 ( .A(
        constructing_unit_Datapath_D_h_4_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n797) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U712 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n797), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n798), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n331) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U711 ( .A(
        constructing_unit_Datapath_D_h_3_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n796) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U710 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n796), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n797), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n332) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U709 ( .A(
        constructing_unit_Datapath_D_h_2_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n795) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U708 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n795), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n796), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n333) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U707 ( .A(
        constructing_unit_Datapath_D_h_1_), .B(
        constructing_unit_Datapath_D_h_11_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n794) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U706 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n794), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n795), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n334) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U705 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n669), .B(
        constructing_unit_Datapath_D_h_0_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n793) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U704 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n793), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n794), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n335) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U703 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n691), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n336) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U702 ( .A(
        constructing_unit_Datapath_n17), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n700) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U701 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n700), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n700), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n792) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U700 ( .A(
        constructing_unit_Datapath_D_h_12_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n791) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U699 ( .A(
        constructing_unit_Datapath_D_h_13_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n697) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U698 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n791), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n697), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n338) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U697 ( .A(
        constructing_unit_Datapath_D_h_11_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n790) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U696 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n790), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n791), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n339) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U695 ( .A(
        constructing_unit_Datapath_D_h_10_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n789) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U694 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n789), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n790), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n340) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U693 ( .A(
        constructing_unit_Datapath_D_h_9_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n788) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U692 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n788), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n789), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n341) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U691 ( .A(
        constructing_unit_Datapath_D_h_8_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n787) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U690 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n787), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n788), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n342) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U689 ( .A(
        constructing_unit_Datapath_D_h_7_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n786) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U688 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n786), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n787), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n343) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U687 ( .A(
        constructing_unit_Datapath_D_h_6_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n785) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U686 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n785), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n786), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n344) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U685 ( .A(
        constructing_unit_Datapath_D_h_5_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n784) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U684 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n784), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n785), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n345) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U683 ( .A(
        constructing_unit_Datapath_D_h_4_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n783) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U682 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n783), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n784), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n346) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U681 ( .A(
        constructing_unit_Datapath_D_h_3_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n782) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U680 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n782), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n783), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n347) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U679 ( .A(
        constructing_unit_Datapath_D_h_2_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n781) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U678 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n781), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n782), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n348) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U677 ( .A(
        constructing_unit_Datapath_D_h_1_), .B(
        constructing_unit_Datapath_D_h_9_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n780) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U676 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n780), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n781), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n349) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U675 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n667), .B(
        constructing_unit_Datapath_D_h_0_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n779) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U674 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n779), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n780), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n350) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U673 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n691), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n351) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U672 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n778), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n778), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n777) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U671 ( .A(
        constructing_unit_Datapath_D_h_12_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n775) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U670 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n775), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n776), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n353) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U669 ( .A(
        constructing_unit_Datapath_D_h_11_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n774) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U668 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n774), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n775), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n354) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U667 ( .A(
        constructing_unit_Datapath_D_h_10_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n773) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U666 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n773), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n774), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n355) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U665 ( .A(
        constructing_unit_Datapath_D_h_9_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n772) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U664 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n772), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n773), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n356) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U663 ( .A(
        constructing_unit_Datapath_D_h_8_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n771) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U662 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n771), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n772), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n357) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U661 ( .A(
        constructing_unit_Datapath_D_h_7_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n770) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U660 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n770), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n771), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n358) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U659 ( .A(
        constructing_unit_Datapath_D_h_6_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n769) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U658 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n769), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n770), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n359) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U657 ( .A(
        constructing_unit_Datapath_D_h_5_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n768) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U656 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n768), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n769), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n360) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U655 ( .A(
        constructing_unit_Datapath_D_h_4_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n767) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U654 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n767), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n768), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n361) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U653 ( .A(
        constructing_unit_Datapath_D_h_3_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n766) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U652 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n766), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n767), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n362) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U651 ( .A(
        constructing_unit_Datapath_D_h_2_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n765) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U650 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n765), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n766), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n363) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U649 ( .A(
        constructing_unit_Datapath_D_h_1_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n764) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U648 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n764), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n765), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n364) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U647 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n665), .B(
        constructing_unit_Datapath_D_h_0_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n762) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U646 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n762), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n764), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n365) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U645 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n691), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n761), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n366) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U644 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n760), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n760), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n759) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U643 ( .A(
        constructing_unit_Datapath_D_h_12_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n757) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U642 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n757), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n758), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n368) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U641 ( .A(
        constructing_unit_Datapath_D_h_11_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n756) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U640 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n756), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n757), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n369) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U639 ( .A(
        constructing_unit_Datapath_D_h_10_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n755) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U638 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n755), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n756), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n370) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U637 ( .A(
        constructing_unit_Datapath_D_h_9_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n754) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U636 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n754), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n755), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n371) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U635 ( .A(
        constructing_unit_Datapath_D_h_8_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n753) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U634 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n753), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n754), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n372) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U633 ( .A(
        constructing_unit_Datapath_D_h_7_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n752) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U632 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n752), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n753), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n373) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U631 ( .A(
        constructing_unit_Datapath_D_h_6_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n751) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U630 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n751), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n752), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n374) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U629 ( .A(
        constructing_unit_Datapath_D_h_5_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n750) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U628 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n750), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n751), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n375) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U627 ( .A(
        constructing_unit_Datapath_D_h_4_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n749) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U626 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n749), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n750), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n376) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U625 ( .A(
        constructing_unit_Datapath_D_h_3_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n748) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U624 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n748), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n749), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n377) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U623 ( .A(
        constructing_unit_Datapath_D_h_2_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n747) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U622 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n747), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n748), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n378) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U621 ( .A(
        constructing_unit_Datapath_D_h_1_), .B(
        constructing_unit_Datapath_D_h_5_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n746) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U620 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n746), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n747), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n379) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U619 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n663), .B(
        constructing_unit_Datapath_D_h_0_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n744) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U618 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n744), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n746), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n380) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U617 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n691), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n743), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n381) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U616 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n742), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n742), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n741) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U615 ( .A(
        constructing_unit_Datapath_D_h_12_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n739) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U614 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n739), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n740), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n383) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U613 ( .A(
        constructing_unit_Datapath_D_h_11_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n738) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U612 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n738), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n739), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n384) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U611 ( .A(
        constructing_unit_Datapath_D_h_10_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n737) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U610 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n737), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n738), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n385) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U609 ( .A(
        constructing_unit_Datapath_D_h_9_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n736) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U608 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n736), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n737), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n386) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U607 ( .A(
        constructing_unit_Datapath_D_h_8_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n735) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U606 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n735), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n736), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n387) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U605 ( .A(
        constructing_unit_Datapath_D_h_7_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n734) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U604 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n734), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n735), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n388) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U603 ( .A(
        constructing_unit_Datapath_D_h_6_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n733) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U602 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n733), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n734), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n389) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U601 ( .A(
        constructing_unit_Datapath_D_h_5_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n732) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U600 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n732), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n733), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n390) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U599 ( .A(
        constructing_unit_Datapath_D_h_4_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n731) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U598 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n731), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n732), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n391) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U597 ( .A(
        constructing_unit_Datapath_D_h_3_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n730) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U596 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n730), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n731), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n392) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U595 ( .A(
        constructing_unit_Datapath_D_h_2_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n729) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U594 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n729), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n730), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n393) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U593 ( .A(
        constructing_unit_Datapath_D_h_1_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n728) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U592 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n728), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n729), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n394) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U591 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n661), .B(
        constructing_unit_Datapath_D_h_0_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n726) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U590 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n726), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n728), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n395) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U589 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n691), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n396) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U588 ( .A(
        constructing_unit_Datapath_n17), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n723) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U587 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n723), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n723), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n724) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U586 ( .A(
        constructing_unit_Datapath_D_h_13_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n722) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U585 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n722), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n723), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n398) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U584 ( .A(
        constructing_unit_Datapath_D_h_12_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n721) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U583 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n721), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n722), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n399) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U582 ( .A(
        constructing_unit_Datapath_D_h_11_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n720) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U581 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n720), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n721), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n400) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U580 ( .A(
        constructing_unit_Datapath_D_h_10_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n719) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U579 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n719), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n720), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n401) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U578 ( .A(
        constructing_unit_Datapath_D_h_9_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n718) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U577 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n718), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n719), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n402) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U576 ( .A(
        constructing_unit_Datapath_D_h_8_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n717) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U575 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n717), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n718), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n403) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U574 ( .A(
        constructing_unit_Datapath_D_h_7_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n716) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U573 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n716), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n717), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n404) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U572 ( .A(
        constructing_unit_Datapath_D_h_6_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n715) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U571 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n715), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n716), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n405) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U570 ( .A(
        constructing_unit_Datapath_D_h_5_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n714) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U569 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n714), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n715), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n406) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U568 ( .A(
        constructing_unit_Datapath_D_h_4_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n713) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U567 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n713), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n714), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n407) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U566 ( .A(
        constructing_unit_Datapath_D_h_3_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n712) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U565 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n712), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n713), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n408) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U564 ( .A(
        constructing_unit_Datapath_D_h_2_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n711) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U563 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n711), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n712), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n409) );
  XNOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U562 ( .A(
        constructing_unit_Datapath_D_h_1_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n710) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U561 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n710), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n711), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n410) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U560 ( .A1(
        constructing_unit_Datapath_D_h_0_), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n710), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n411) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U559 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n705), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n708), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n70) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U558 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n701), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n704), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n80) );
  OAI22_X1 constructing_unit_Datapath_L_squarer_mult_13_U557 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n697), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n700), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n94) );
  NOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U556 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n691), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_D_h_sq_tmp[0]) );
  XOR2_X1 constructing_unit_Datapath_L_squarer_mult_13_U555 ( .A(
        constructing_unit_Datapath_n17), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n674), .Z(
        constructing_unit_Datapath_L_squarer_mult_13_n696) );
  NAND2_X1 constructing_unit_Datapath_L_squarer_mult_13_U554 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n696), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n689), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n693) );
  AOI222_X1 constructing_unit_Datapath_L_squarer_mult_13_U553 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n38), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n68), .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n38), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n67), .C1(
        constructing_unit_Datapath_L_squarer_mult_13_n67), .C2(
        constructing_unit_Datapath_L_squarer_mult_13_n68), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n695) );
  AND2_X1 constructing_unit_Datapath_L_squarer_mult_13_U552 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n693), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n675), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n694) );
  AOI221_X1 constructing_unit_Datapath_L_squarer_mult_13_U551 ( .B1(
        constructing_unit_Datapath_L_squarer_mult_13_n66), .B2(
        constructing_unit_Datapath_L_squarer_mult_13_n693), .C1(
        constructing_unit_Datapath_L_squarer_mult_13_n66), .C2(
        constructing_unit_Datapath_L_squarer_mult_13_n675), .A(
        constructing_unit_Datapath_L_squarer_mult_13_n694), .ZN(
        constructing_unit_Datapath_L_squarer_product_29_) );
  INV_X2 constructing_unit_Datapath_L_squarer_mult_13_U550 ( .A(
        constructing_unit_Datapath_D_h_0_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n692) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U549 ( .A(
        constructing_unit_Datapath_D_h_13_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n672) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U548 ( .A(
        constructing_unit_Datapath_D_h_11_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n670) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U547 ( .A(
        constructing_unit_Datapath_D_h_9_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n668) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U546 ( .A(
        constructing_unit_Datapath_D_h_7_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n666) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U545 ( .A(
        constructing_unit_Datapath_D_h_5_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n664) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U544 ( .A(
        constructing_unit_Datapath_D_h_3_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n662) );
  XOR2_X2 constructing_unit_Datapath_L_squarer_mult_13_U543 ( .A(
        constructing_unit_Datapath_D_h_6_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n664), .Z(
        constructing_unit_Datapath_L_squarer_mult_13_n761) );
  XOR2_X2 constructing_unit_Datapath_L_squarer_mult_13_U542 ( .A(
        constructing_unit_Datapath_D_h_4_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n662), .Z(
        constructing_unit_Datapath_L_squarer_mult_13_n743) );
  XOR2_X2 constructing_unit_Datapath_L_squarer_mult_13_U541 ( .A(
        constructing_unit_Datapath_D_h_2_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n660), .Z(
        constructing_unit_Datapath_L_squarer_mult_13_n725) );
  XOR2_X2 constructing_unit_Datapath_L_squarer_mult_13_U540 ( .A(
        constructing_unit_Datapath_D_h_12_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n670), .Z(
        constructing_unit_Datapath_L_squarer_mult_13_n707) );
  XOR2_X2 constructing_unit_Datapath_L_squarer_mult_13_U539 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n674), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n672), .Z(
        constructing_unit_Datapath_L_squarer_mult_13_n821) );
  XOR2_X2 constructing_unit_Datapath_L_squarer_mult_13_U538 ( .A(
        constructing_unit_Datapath_D_h_10_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n668), .Z(
        constructing_unit_Datapath_L_squarer_mult_13_n703) );
  XOR2_X2 constructing_unit_Datapath_L_squarer_mult_13_U537 ( .A(
        constructing_unit_Datapath_D_h_8_), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n666), .Z(
        constructing_unit_Datapath_L_squarer_mult_13_n699) );
  NAND2_X2 constructing_unit_Datapath_L_squarer_mult_13_U536 ( .A1(
        constructing_unit_Datapath_L_squarer_mult_13_n725), .A2(
        constructing_unit_Datapath_L_squarer_mult_13_n846), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n727) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U535 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n70), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n682) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U534 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n759), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n686) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U533 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n741), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n684) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U532 ( .A(
        constructing_unit_Datapath_D_h_1_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n660) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U531 ( .A(
        constructing_unit_Datapath_D_h_0_), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n691) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U530 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n695), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n675) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U529 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n820), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n681) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U528 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n806), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n679) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U527 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n777), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n688) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U526 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n112), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n687) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U525 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n792), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n677) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U524 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n80), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n680) );
  BUF_X1 constructing_unit_Datapath_L_squarer_mult_13_U523 ( .A(
        constructing_unit_Datapath_n17), .Z(
        constructing_unit_Datapath_L_squarer_mult_13_n673) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U522 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n844), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n690) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U521 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n134), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n685) );
  BUF_X1 constructing_unit_Datapath_L_squarer_mult_13_U520 ( .A(
        constructing_unit_Datapath_n17), .Z(
        constructing_unit_Datapath_L_squarer_mult_13_n674) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U519 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n160), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n683) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U518 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n724), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n676) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U517 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n660), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n659) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U516 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n662), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n661) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U515 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n666), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n665) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U514 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n664), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n663) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U513 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n668), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n667) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U512 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n672), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n671) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U511 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n670), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n669) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U510 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n94), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n678) );
  INV_X1 constructing_unit_Datapath_L_squarer_mult_13_U509 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n821), .ZN(
        constructing_unit_Datapath_L_squarer_mult_13_n689) );
  HA_X1 constructing_unit_Datapath_L_squarer_mult_13_U163 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n395), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n409), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n258), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n259) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U162 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n408), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n381), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n394), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n256), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n257) );
  HA_X1 constructing_unit_Datapath_L_squarer_mult_13_U161 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n289), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n380), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n254), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n255) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U160 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n393), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n407), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n255), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n252), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n253) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U159 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n406), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n366), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n392), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n250), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n251) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U158 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n254), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n379), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n251), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n248), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n249) );
  HA_X1 constructing_unit_Datapath_L_squarer_mult_13_U157 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n288), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n365), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n246), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n247) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U156 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n378), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n405), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n391), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n244), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n245) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U155 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n250), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n247), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n245), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n242), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n243) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U154 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n377), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n351), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n404), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n240), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n241) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U153 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n364), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n390), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n246), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n238), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n239) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U152 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n241), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n244), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n239), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n236), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n237) );
  HA_X1 constructing_unit_Datapath_L_squarer_mult_13_U151 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n287), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n350), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n234), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n235) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U150 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n363), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n376), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n389), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n232), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n233) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U149 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n235), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n403), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n240), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n230), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n231) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U148 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n233), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n238), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n231), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n228), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n229) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U147 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n362), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n336), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n402), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n226), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n227) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U146 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n349), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n388), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n375), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n224), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n225) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U145 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n232), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n234), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n227), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n222), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n223) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U144 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n230), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n225), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n223), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n220), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n221) );
  HA_X1 constructing_unit_Datapath_L_squarer_mult_13_U143 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n286), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n335), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n218), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n219) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U142 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n348), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n374), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n401), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n216), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n217) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U141 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n361), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n387), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n219), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n214), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n215) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U140 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n224), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n226), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n217), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n212), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n213) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U139 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n222), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n215), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n213), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n210), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n211) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U138 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n347), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n321), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n400), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n208), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n209) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U137 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n334), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n386), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n360), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n206), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n207) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U136 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n218), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n373), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n216), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n204), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n205) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U135 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n207), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n209), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n214), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n202), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n203) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U134 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n205), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n212), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n203), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n200), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n201) );
  HA_X1 constructing_unit_Datapath_L_squarer_mult_13_U133 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n285), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n320), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n198), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n199) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U132 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n399), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n359), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n385), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n196), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n197) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U131 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n333), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n372), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n346), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n194), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n195) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U130 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n208), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n199), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n206), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n192), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n193) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U129 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n197), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n195), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n204), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n190), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n191) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U128 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n202), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n193), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n191), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n188), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n189) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U127 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n332), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n306), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n398), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n186), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n187) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U126 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n319), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n384), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n345), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n184), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n185) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U125 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n358), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n371), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n198), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n182), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n183) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U124 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n194), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n196), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n187), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n180), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n181) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U123 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n183), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n185), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n192), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n178), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n179) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U122 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n181), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n190), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n179), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n176), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n177) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U119 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n284), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n357), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n676), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n172), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n173) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U118 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n383), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n331), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n344), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n170), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n171) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U117 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n175), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n370), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n186), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n168), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n169) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U116 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n182), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n184), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n171), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n166), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n167) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U115 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n180), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n173), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n169), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n164), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n165) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U114 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n167), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n178), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n165), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n162), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n163) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U112 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n369), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n330), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n304), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n158), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n159) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U111 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n317), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n356), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n343), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n156), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n157) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U110 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n174), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n683), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n172), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n154), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n155) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U109 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n157), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n170), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n159), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n152), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n153) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U108 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n166), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n168), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n155), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n150), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n151) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U107 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n164), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n153), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n151), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n148), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n149) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U106 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n160), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n303), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n684), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n146), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n147) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U105 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n316), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n368), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n355), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n144), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n145) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U104 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n329), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n342), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n158), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n142), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n143) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U103 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n145), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n156), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n147), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n140), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n141) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U102 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n143), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n154), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n152), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n138), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n139) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U101 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n150), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n141), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n139), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n136), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n137) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U99 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n354), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n328), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n341), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n132), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n133) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U98 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n302), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n315), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n685), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n130), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n131) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U97 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n144), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n146), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n133), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n128), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n129) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U96 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n142), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n131), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n140), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n126), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n127) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U95 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n138), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n129), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n127), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n124), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n125) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U94 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n134), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n301), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n686), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n122), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n123) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U93 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n314), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n353), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n327), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n120), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n121) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U92 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n132), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n340), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n130), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n118), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n119) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U91 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n123), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n121), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n128), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n116), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n117) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U90 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n126), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n119), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n117), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n114), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n115) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U88 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n339), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n313), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n300), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n110), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n111) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U87 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n687), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n326), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n122), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n108), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n109) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U86 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n111), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n120), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n118), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n106), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n107) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U85 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n116), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n109), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n107), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n104), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n105) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U84 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n338), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n299), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n688), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n102), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n103) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U83 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n312), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n112), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n325), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n100), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n101) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U82 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n101), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n110), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n103), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n98), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n99) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U81 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n106), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n108), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n99), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n96), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n97) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U79 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n298), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n311), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n324), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n92), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n93) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U78 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n102), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n678), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n100), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n90), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n91) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U77 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n91), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n93), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n98), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n88), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n89) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U76 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n310), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n297), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n677), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n86), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n87) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U75 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n94), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n323), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n92), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n84), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n85) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U74 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n90), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n87), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n85), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n82), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n83) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U72 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n296), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n309), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n680), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n78), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n79) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U71 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n79), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n86), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n84), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n76), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n77) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U70 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n308), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n80), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n679), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n74), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n75) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U69 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n78), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n295), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n75), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n72), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n73) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U67 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n682), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n294), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n74), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n68), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n69) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U66 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n293), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n70), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n681), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n66), .S(
        constructing_unit_Datapath_L_squarer_mult_13_n67) );
  HA_X1 constructing_unit_Datapath_L_squarer_mult_13_U64 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n411), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n291), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n63), .S(
        constructing_unit_Datapath_D_h_sq_tmp[1]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U63 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n410), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n396), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n63), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n62), .S(
        constructing_unit_Datapath_D_h_sq_tmp[2]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U62 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n259), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n290), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n62), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n61), .S(
        constructing_unit_Datapath_D_h_sq_tmp[3]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U61 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n257), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n258), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n61), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n60), .S(
        constructing_unit_Datapath_D_h_sq_tmp[4]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U60 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n253), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n256), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n60), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n59), .S(
        constructing_unit_Datapath_D_h_sq_tmp[5]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U59 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n249), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n252), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n59), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n58), .S(
        constructing_unit_Datapath_D_h_sq_tmp[6]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U58 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n243), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n248), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n58), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n57), .S(
        constructing_unit_Datapath_D_h_sq_tmp[7]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U57 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n237), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n242), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n57), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n56), .S(
        constructing_unit_Datapath_D_h_sq_tmp[8]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U56 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n229), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n236), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n56), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n55), .S(
        constructing_unit_Datapath_D_h_sq_tmp[9]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U55 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n221), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n228), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n55), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n54), .S(
        constructing_unit_Datapath_D_h_sq_tmp[10]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U54 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n211), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n220), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n54), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n53), .S(
        constructing_unit_Datapath_D_h_sq_tmp[11]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U53 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n201), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n210), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n53), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n52), .S(
        constructing_unit_Datapath_D_h_sq_tmp[12]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U52 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n189), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n200), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n52), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n51), .S(
        constructing_unit_Datapath_D_h_sq_tmp[13]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U51 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n177), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n188), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n51), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n50), .S(
        constructing_unit_Datapath_D_h_sq_tmp[14]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U50 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n163), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n176), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n50), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n49), .S(
        constructing_unit_Datapath_D_h_sq_tmp[15]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U49 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n149), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n162), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n49), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n48), .S(
        constructing_unit_Datapath_D_h_sq_tmp[16]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U48 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n137), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n148), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n48), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n47), .S(
        constructing_unit_Datapath_D_h_sq_tmp[17]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U47 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n125), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n136), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n47), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n46), .S(
        constructing_unit_Datapath_D_h_sq_tmp[18]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U46 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n115), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n124), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n46), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n45), .S(
        constructing_unit_Datapath_D_h_sq_tmp[19]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U45 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n105), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n114), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n45), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n44), .S(
        constructing_unit_Datapath_D_h_sq_tmp[20]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U44 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n97), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n104), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n44), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n43), .S(
        constructing_unit_Datapath_D_h_sq_tmp[21]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U43 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n89), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n96), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n43), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n42), .S(
        constructing_unit_Datapath_D_h_sq_tmp[22]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U42 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n83), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n88), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n42), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n41), .S(
        constructing_unit_Datapath_D_h_sq_tmp[23]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U41 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n77), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n82), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n41), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n40), .S(
        constructing_unit_Datapath_D_h_sq_tmp[24]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U40 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n73), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n76), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n40), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n39), .S(
        constructing_unit_Datapath_D_h_sq_tmp[25]) );
  FA_X1 constructing_unit_Datapath_L_squarer_mult_13_U39 ( .A(
        constructing_unit_Datapath_L_squarer_mult_13_n69), .B(
        constructing_unit_Datapath_L_squarer_mult_13_n72), .CI(
        constructing_unit_Datapath_L_squarer_mult_13_n39), .CO(
        constructing_unit_Datapath_L_squarer_mult_13_n38), .S(
        constructing_unit_Datapath_D_h_sq_tmp[26]) );
  INV_X1 constructing_unit_Datapath_R_sub1_sub_19_U14 ( .A(
        constructing_unit_Datapath_MV0_int_h_1__10_), .ZN(
        constructing_unit_Datapath_R_sub1_sub_19_n2) );
  XNOR2_X1 constructing_unit_Datapath_R_sub1_sub_19_U13 ( .A(
        constructing_unit_Datapath_R_sub1_sub_19_n12), .B(
        constructing_unit_Datapath_MV1_int_h_1__0_), .ZN(
        constructing_unit_Datapath_mv1h_mv0h_int[0]) );
  INV_X1 constructing_unit_Datapath_R_sub1_sub_19_U12 ( .A(
        constructing_unit_Datapath_MV0_int_h_1__0_), .ZN(
        constructing_unit_Datapath_R_sub1_sub_19_n12) );
  INV_X1 constructing_unit_Datapath_R_sub1_sub_19_U11 ( .A(
        constructing_unit_Datapath_MV0_int_h_1__9_), .ZN(
        constructing_unit_Datapath_R_sub1_sub_19_n3) );
  INV_X1 constructing_unit_Datapath_R_sub1_sub_19_U10 ( .A(
        constructing_unit_Datapath_MV0_int_h_1__8_), .ZN(
        constructing_unit_Datapath_R_sub1_sub_19_n4) );
  INV_X1 constructing_unit_Datapath_R_sub1_sub_19_U9 ( .A(
        constructing_unit_Datapath_MV0_int_h_1__7_), .ZN(
        constructing_unit_Datapath_R_sub1_sub_19_n5) );
  INV_X1 constructing_unit_Datapath_R_sub1_sub_19_U8 ( .A(
        constructing_unit_Datapath_MV0_int_h_1__6_), .ZN(
        constructing_unit_Datapath_R_sub1_sub_19_n6) );
  INV_X1 constructing_unit_Datapath_R_sub1_sub_19_U7 ( .A(
        constructing_unit_Datapath_MV0_int_h_1__5_), .ZN(
        constructing_unit_Datapath_R_sub1_sub_19_n7) );
  INV_X1 constructing_unit_Datapath_R_sub1_sub_19_U6 ( .A(
        constructing_unit_Datapath_MV0_int_h_1__4_), .ZN(
        constructing_unit_Datapath_R_sub1_sub_19_n8) );
  INV_X1 constructing_unit_Datapath_R_sub1_sub_19_U5 ( .A(
        constructing_unit_Datapath_MV0_int_h_1__3_), .ZN(
        constructing_unit_Datapath_R_sub1_sub_19_n9) );
  INV_X1 constructing_unit_Datapath_R_sub1_sub_19_U4 ( .A(
        constructing_unit_Datapath_MV0_int_h_1__2_), .ZN(
        constructing_unit_Datapath_R_sub1_sub_19_n10) );
  INV_X1 constructing_unit_Datapath_R_sub1_sub_19_U3 ( .A(
        constructing_unit_Datapath_MV1_int_h_1__0_), .ZN(
        constructing_unit_Datapath_R_sub1_sub_19_n1) );
  NAND2_X1 constructing_unit_Datapath_R_sub1_sub_19_U2 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__0_), .A2(
        constructing_unit_Datapath_R_sub1_sub_19_n1), .ZN(
        constructing_unit_Datapath_R_sub1_sub_19_carry[1]) );
  INV_X1 constructing_unit_Datapath_R_sub1_sub_19_U1 ( .A(
        constructing_unit_Datapath_MV0_int_h_1__1_), .ZN(
        constructing_unit_Datapath_R_sub1_sub_19_n11) );
  FA_X1 constructing_unit_Datapath_R_sub1_sub_19_U2_1 ( .A(
        constructing_unit_Datapath_MV1_int_h_1__1_), .B(
        constructing_unit_Datapath_R_sub1_sub_19_n11), .CI(
        constructing_unit_Datapath_R_sub1_sub_19_carry[1]), .CO(
        constructing_unit_Datapath_R_sub1_sub_19_carry[2]), .S(
        constructing_unit_Datapath_mv1h_mv0h_int[1]) );
  FA_X1 constructing_unit_Datapath_R_sub1_sub_19_U2_2 ( .A(
        constructing_unit_Datapath_MV1_int_h_1__2_), .B(
        constructing_unit_Datapath_R_sub1_sub_19_n10), .CI(
        constructing_unit_Datapath_R_sub1_sub_19_carry[2]), .CO(
        constructing_unit_Datapath_R_sub1_sub_19_carry[3]), .S(
        constructing_unit_Datapath_mv1h_mv0h_int[2]) );
  FA_X1 constructing_unit_Datapath_R_sub1_sub_19_U2_3 ( .A(
        constructing_unit_Datapath_MV1_int_h_1__3_), .B(
        constructing_unit_Datapath_R_sub1_sub_19_n9), .CI(
        constructing_unit_Datapath_R_sub1_sub_19_carry[3]), .CO(
        constructing_unit_Datapath_R_sub1_sub_19_carry[4]), .S(
        constructing_unit_Datapath_mv1h_mv0h_int[3]) );
  FA_X1 constructing_unit_Datapath_R_sub1_sub_19_U2_4 ( .A(
        constructing_unit_Datapath_MV1_int_h_1__4_), .B(
        constructing_unit_Datapath_R_sub1_sub_19_n8), .CI(
        constructing_unit_Datapath_R_sub1_sub_19_carry[4]), .CO(
        constructing_unit_Datapath_R_sub1_sub_19_carry[5]), .S(
        constructing_unit_Datapath_mv1h_mv0h_int[4]) );
  FA_X1 constructing_unit_Datapath_R_sub1_sub_19_U2_5 ( .A(
        constructing_unit_Datapath_MV1_int_h_1__5_), .B(
        constructing_unit_Datapath_R_sub1_sub_19_n7), .CI(
        constructing_unit_Datapath_R_sub1_sub_19_carry[5]), .CO(
        constructing_unit_Datapath_R_sub1_sub_19_carry[6]), .S(
        constructing_unit_Datapath_mv1h_mv0h_int[5]) );
  FA_X1 constructing_unit_Datapath_R_sub1_sub_19_U2_6 ( .A(
        constructing_unit_Datapath_MV1_int_h_1__6_), .B(
        constructing_unit_Datapath_R_sub1_sub_19_n6), .CI(
        constructing_unit_Datapath_R_sub1_sub_19_carry[6]), .CO(
        constructing_unit_Datapath_R_sub1_sub_19_carry[7]), .S(
        constructing_unit_Datapath_mv1h_mv0h_int[6]) );
  FA_X1 constructing_unit_Datapath_R_sub1_sub_19_U2_7 ( .A(
        constructing_unit_Datapath_MV1_int_h_1__7_), .B(
        constructing_unit_Datapath_R_sub1_sub_19_n5), .CI(
        constructing_unit_Datapath_R_sub1_sub_19_carry[7]), .CO(
        constructing_unit_Datapath_R_sub1_sub_19_carry[8]), .S(
        constructing_unit_Datapath_mv1h_mv0h_int[7]) );
  FA_X1 constructing_unit_Datapath_R_sub1_sub_19_U2_8 ( .A(
        constructing_unit_Datapath_MV1_int_h_1__8_), .B(
        constructing_unit_Datapath_R_sub1_sub_19_n4), .CI(
        constructing_unit_Datapath_R_sub1_sub_19_carry[8]), .CO(
        constructing_unit_Datapath_R_sub1_sub_19_carry[9]), .S(
        constructing_unit_Datapath_mv1h_mv0h_int[8]) );
  FA_X1 constructing_unit_Datapath_R_sub1_sub_19_U2_9 ( .A(
        constructing_unit_Datapath_MV1_int_h_1__9_), .B(
        constructing_unit_Datapath_R_sub1_sub_19_n3), .CI(
        constructing_unit_Datapath_R_sub1_sub_19_carry[9]), .CO(
        constructing_unit_Datapath_R_sub1_sub_19_carry[10]), .S(
        constructing_unit_Datapath_mv1h_mv0h_int[9]) );
  FA_X1 constructing_unit_Datapath_R_sub1_sub_19_U2_10 ( .A(
        constructing_unit_Datapath_MV1_int_h_1__10_), .B(
        constructing_unit_Datapath_R_sub1_sub_19_n2), .CI(
        constructing_unit_Datapath_R_sub1_sub_19_carry[10]), .CO(
        constructing_unit_Datapath_R_sub1_sub_19_carry[11]), .S(
        constructing_unit_Datapath_mv1h_mv0h_int[10]) );
  FA_X1 constructing_unit_Datapath_R_sub1_sub_19_U2_11 ( .A(
        constructing_unit_Datapath_MV1_int_h_1__10_), .B(
        constructing_unit_Datapath_R_sub1_sub_19_n2), .CI(
        constructing_unit_Datapath_R_sub1_sub_19_carry[11]), .S(
        constructing_unit_Datapath_mv1h_mv0h_int[11]) );
  INV_X1 constructing_unit_Datapath_mv1h_mv0h_REG_0_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_mv1h_mv0h_REG_0_n1) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_0_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[0]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[12]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_0_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[1]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[13]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_0_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[2]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[14]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_0_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[3]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[15]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_0_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[4]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[16]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_0_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[5]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[17]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_0_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[6]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[18]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_0_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[7]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[19]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_0_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[8]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[20]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_0_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[9]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[21]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_0_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[10]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[22]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_0_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[11]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_0_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[23]) );
  INV_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_2_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_2_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[12]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[24]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_2_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[13]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[25]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_2_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[14]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[26]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_2_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[15]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[27]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_2_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[16]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[28]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_2_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[17]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[29]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_2_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[18]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[30]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_2_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[19]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[31]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_2_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[20]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[32]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_2_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[21]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[33]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_2_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[22]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[34]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_2_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[23]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_2_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[35]) );
  INV_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_3_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_3_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[24]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[36]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_3_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[25]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[37]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_3_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[26]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[38]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_3_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[27]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[39]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_3_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[28]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[40]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_3_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[29]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[41]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_3_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[30]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[42]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_3_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[31]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[43]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_3_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[32]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[44]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_3_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[33]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[45]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_3_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[34]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[46]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_3_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[35]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_3_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[47]) );
  INV_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_4_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_4_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[36]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[48]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_4_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[37]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[49]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_4_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[38]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[50]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_4_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[39]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[51]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_4_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[40]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[52]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_4_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[41]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[53]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_4_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[42]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[54]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_4_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[43]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[55]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_4_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[44]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[56]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_4_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[45]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[57]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_4_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[46]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[58]) );
  DFFR_X1 constructing_unit_Datapath_mv1h_mv0h_REG_X_4_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_mv1h_mv0h_int[47]), .CK(clk), .RN(
        constructing_unit_Datapath_mv1h_mv0h_REG_X_4_n1), .Q(
        constructing_unit_Datapath_mv1h_mv0h_int[59]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U33 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[13]), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[13]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n35) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U32 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n35), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[13]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U31 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[12]), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[13]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n34) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U30 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n34), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[12]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U29 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[11]), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[13]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n33) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U28 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n33), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[11]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U27 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[10]), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[10]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n32) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U26 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n32), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[10]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U25 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[8]), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[8]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n43) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U24 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n43), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[8]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U23 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[7]), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[7]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n42) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U22 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n42), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[7]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U21 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[6]), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[6]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n41) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U20 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n41), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[6]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U19 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[5]), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[5]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n40) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U18 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n40), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[5]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U17 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[4]), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[4]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n39) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U16 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n39), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[4]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U15 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[3]), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[3]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n38) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U14 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n38), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[3]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U13 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[2]), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[2]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n37) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U12 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n37), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[2]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U11 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[1]), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[1]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n36) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U10 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n36), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[1]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U9 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[0]), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[0]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n31) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U8 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n31), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[0]) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_U7 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .A2(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[9]), .B1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[9]), .B2(
        constructing_unit_Datapath_R_LR_SH2_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n44) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U6 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n44), .ZN(
        constructing_unit_Datapath_diff_mult_h_int[9]) );
  OR2_X1 constructing_unit_Datapath_R_LR_SH2_U5 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_shift_amt_int_0_), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_amt_int_1_), .ZN(
        constructing_unit_Datapath_R_LR_SH2_SH_en) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U4 ( .A(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_1_), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n15) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_U3 ( .A(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_), .ZN(
        constructing_unit_Datapath_R_LR_SH2_n16) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_FF_X_1_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_R_LR_SH2_FF_X_1_n1) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_FF_X_1_Q_int_reg ( .D(
        constructing_unit_Datapath_SH_cmd_int_2_), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_FF_X_1_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_1_) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_FF_X_2_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_R_LR_SH2_FF_X_2_n1) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_FF_X_2_Q_int_reg ( .D(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_1_), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_FF_X_2_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_2_) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_FF_X_3_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_R_LR_SH2_FF_X_3_n1) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_FF_X_3_Q_int_reg ( .D(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_2_), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_FF_X_3_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_3_) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_shift_amt_sample_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_R_LR_SH2_shift_amt_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_shift_amt_sample_Q_int_reg_0_ ( 
        .D(constructing_unit_Datapath_SH_cmd_int_0_), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_shift_amt_sample_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_shift_amt_int_0_) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_shift_amt_sample_Q_int_reg_1_ ( 
        .D(constructing_unit_Datapath_SH_cmd_int_1_), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_shift_amt_sample_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_shift_amt_int_1_) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_SH_en2_sampling_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_R_LR_SH2_SH_en2_sampling_n1) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_SH_en2_sampling_Q_int_reg ( .D(
        constructing_unit_Datapath_R_LR_SH2_shift_amt_int_1_), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_SH_en2_sampling_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_SH_en2) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U40 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n1) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U39 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_n15), .A2(
        constructing_unit_Datapath_mv1h_mv0h_int[59]), .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n16), .B2(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[11]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n52) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U38 ( .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n52), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n2) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U37 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[58]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n5) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U36 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[57]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n6) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U35 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[56]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n7) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U34 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[55]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n8) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U33 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[54]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n9) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U32 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[53]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n10) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U31 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[52]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n11) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U30 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[51]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n12) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U29 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[50]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n13) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U28 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[49]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n14) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U27 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[10]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n53) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U26 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[59]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n4) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U25 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n5), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n4), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n53), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n41) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U24 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[9]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n54) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U23 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n6), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n5), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n54), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n42) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U22 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[8]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n55) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U21 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n7), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n6), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n55), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n43) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U20 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[7]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n56) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U19 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n8), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n7), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n56), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n44) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U18 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[6]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n57) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U17 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n9), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n8), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n57), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n45) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U16 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[5]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n58) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U15 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n10), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n9), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n58), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n46) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U14 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[4]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n59) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U13 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n11), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n10), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n59), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n47) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U12 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[3]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n60) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U11 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n12), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n11), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n60), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n48) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U10 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[2]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n61) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U9 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n13), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n12), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n61), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n49) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U8 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[1]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n62) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U7 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n14), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n13), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n62), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n50) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U6 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[48]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n15) );
  OAI222_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U5 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n65), .A2(
        constructing_unit_Datapath_R_LR_SH2_n15), .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n15), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n64), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n14), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n63), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n51) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U4 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_SH_en), .A2(
        constructing_unit_Datapath_R_LR_SH2_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n63) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U3 ( .A(
        constructing_unit_Datapath_R_LR_SH2_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n16) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_U2 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_n15), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n63), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n64) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_SH_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_first_n51), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[0]), .QN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n65) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_SH_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_first_n50), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[1]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_SH_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_first_n49), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[2]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_SH_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_first_n48), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[3]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_SH_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_first_n47), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[4]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_SH_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_first_n46), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[5]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_SH_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_first_n45), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[6]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_SH_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_first_n44), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[7]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_SH_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_first_n43), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[8]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_SH_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_first_n42), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[9]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_SH_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_first_n41), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[10]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_first_SH_out_int_reg_11_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_first_n2), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[11]) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U40 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n1) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U39 ( .A(1'b1), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n16) );
  AOI22_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U38 ( .A1(1'b1), 
        .A2(constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[11]), .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n16), .B2(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[13]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n52) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U37 ( .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n52), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n4) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U36 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[10]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n5) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U35 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[9]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n6) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U34 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[8]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n7) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U33 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[7]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n8) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U32 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[6]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n9) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U31 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[5]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n10) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U30 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[4]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n11) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U29 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[3]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n12) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U28 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[2]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n13) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U27 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[1]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n14) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U26 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[11]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n2) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U25 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[10]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n53) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U24 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n5), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n2), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n53), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n41) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U23 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[9]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n54) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U22 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n6), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n5), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n54), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n42) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U21 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[8]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n55) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U20 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n7), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n6), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n55), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n43) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U19 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[7]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n56) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U18 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n8), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n7), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n56), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n44) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U17 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[6]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n57) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U16 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n9), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n8), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n57), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n45) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U15 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[5]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n58) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U14 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n10), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n9), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n58), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n46) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U13 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[4]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n59) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U12 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n11), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n10), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n59), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n47) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U11 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[3]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n60) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U10 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n12), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n11), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n60), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n48) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U9 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[2]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n61) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U8 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n13), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n12), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n61), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n49) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U7 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[1]), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n62) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U6 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n64), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n14), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n63), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n13), .A(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n62), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n50) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U5 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1R[0]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n15) );
  OAI222_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U4 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n65), .A2(1'b1), .B1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n15), .B2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n64), .C1(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n14), .C2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n63), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n51) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U3 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_SH_en2), .A2(1'b1), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n63) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_U2 ( .A1(1'b1), .A2(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n63), .ZN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n64) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_SH_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_second_n51), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[0]), .QN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n65) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_SH_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_second_n50), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[1]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_SH_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_second_n49), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[2]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_SH_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_second_n48), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[3]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_SH_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_second_n47), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[4]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_SH_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_second_n46), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[5]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_SH_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_second_n45), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[6]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_SH_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_second_n44), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[7]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_SH_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_second_n43), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[8]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_SH_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_second_n42), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[9]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_SH_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_second_n41), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[10]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_RSH_second_SH_out_int_reg_11_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_RSH_second_n4), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_RSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2R_ext[13]) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U42 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U41 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[58]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n4) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U40 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[57]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n5) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U39 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[56]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n6) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U38 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[55]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n7) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U37 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[54]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n8) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U36 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[53]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n9) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U35 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[52]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n10) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U34 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[51]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n11) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U33 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[50]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n12) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U32 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[49]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n13) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U31 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[48]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n14) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U30 ( .A(
        constructing_unit_Datapath_mv1h_mv0h_int[59]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n3) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U29 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[0]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n68) );
  OAI21_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U28 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n69), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n14), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n68), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n55) );
  OAI22_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U27 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n3), .B1(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_1_), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n70), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n43) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U26 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[1]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n66) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U25 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n14), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n67), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n69), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n13), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n66), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n54) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U24 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[11]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n56) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U23 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n67), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n4), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n69), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n3), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n56), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n44) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U22 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[10]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n57) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U21 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n67), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n5), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n69), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n4), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n57), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n45) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U20 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[9]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n58) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U19 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n67), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n6), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n69), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n5), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n58), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n46) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U18 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[8]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n59) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U17 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n67), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n7), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n69), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n6), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n59), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n47) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U16 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[7]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n60) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U15 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n67), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n8), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n69), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n7), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n60), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n48) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U14 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[6]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n61) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U13 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n67), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n9), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n69), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n8), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n61), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n49) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U12 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[5]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n62) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U11 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n67), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n10), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n69), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n9), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n62), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n50) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U10 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[4]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n63) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U9 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n67), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n11), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n69), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n10), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n63), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n51) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U8 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[3]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n64) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U7 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n67), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n12), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n69), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n11), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n64), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n52) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U6 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[2]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n65) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U5 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n67), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n13), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n69), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n12), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n65), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n53) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U4 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_1_), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n67), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n69) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U3 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_SH_en), .A2(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_1_), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n67) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_U2 ( .A(
        constructing_unit_Datapath_R_LR_SH2_shift_dir_int_1_), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n15) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_SH_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_first_n55), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[0]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_SH_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_first_n54), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[1]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_SH_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_first_n53), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[2]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_SH_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_first_n52), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[3]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_SH_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_first_n51), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[4]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_SH_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_first_n50), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[5]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_SH_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_first_n49), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[6]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_SH_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_first_n48), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[7]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_SH_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_first_n47), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[8]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_SH_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_first_n46), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[9]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_SH_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_first_n45), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[10]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_SH_out_int_reg_11_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_first_n44), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[11]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_first_SH_out_int_reg_12_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_first_n43), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[12]), .QN(
        constructing_unit_Datapath_R_LR_SH2_LSH_first_n70) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U45 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U44 ( .A(1'b1), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U43 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[12]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n3) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U42 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[11]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n4) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U41 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[10]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n5) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U40 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[9]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n6) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U39 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[8]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n7) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U38 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[7]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n8) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U37 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[6]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n9) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U36 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[5]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n10) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U35 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[4]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n11) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U34 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[3]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n12) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U33 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[2]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n13) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U32 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[1]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n14) );
  INV_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U31 ( .A(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d1L[0]), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n15) );
  OAI22_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U30 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n3), .B1(1'b1), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n75), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n46) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U29 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[0]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n73) );
  OAI21_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U28 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n15), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n73), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n59) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U27 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[1]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n71) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U26 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n15), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n14), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n71), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n58) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U25 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[12]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n60) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U24 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n4), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n3), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n60), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n47) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U23 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[11]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n61) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U22 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n5), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n4), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n61), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n48) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U21 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[10]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n62) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U20 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n6), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n5), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n62), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n49) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U19 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[9]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n63) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U18 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n7), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n6), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n63), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n50) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U17 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[8]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n64) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U16 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n8), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n7), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n64), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n51) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U15 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[7]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n65) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U14 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n9), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n8), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n65), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n52) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U13 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[6]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n66) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U12 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n10), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n9), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n66), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n53) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U11 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[5]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n67) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U10 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n11), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n10), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n67), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n54) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U9 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[4]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n68) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U8 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n12), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n11), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n68), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n55) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U7 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[3]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n69) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U6 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n13), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n12), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n69), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n56) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U5 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[2]), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n16), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n70) );
  OAI221_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U4 ( .B1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72), .B2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n14), .C1(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74), .C2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n13), .A(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n70), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n57) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U3 ( .A1(1'b1), .A2(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n74) );
  NAND2_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_U2 ( .A1(
        constructing_unit_Datapath_R_LR_SH2_SH_en2), .A2(1'b1), .ZN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n72) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n59), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[0]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n58), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[1]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n57), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[2]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n56), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[3]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n55), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[4]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n54), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[5]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n53), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[6]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n52), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[7]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n51), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[8]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n50), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[9]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n49), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[10]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_11_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n48), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[11]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_12_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n47), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[12]) );
  DFFR_X1 constructing_unit_Datapath_R_LR_SH2_LSH_second_SH_out_int_reg_13_ ( 
        .D(constructing_unit_Datapath_R_LR_SH2_LSH_second_n46), .CK(clk), .RN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n1), .Q(
        constructing_unit_Datapath_R_LR_SH2_MV1_MV0_d2L[13]), .QN(
        constructing_unit_Datapath_R_LR_SH2_LSH_second_n75) );
  INV_X1 constructing_unit_Datapath_diff_mult_h_int_samp_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[0]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[14]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[1]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[15]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[2]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[16]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[3]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[17]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[4]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[18]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[5]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[19]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[6]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[20]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[7]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[21]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[8]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[22]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[9]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[23]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[10]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[24]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[11]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[25]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[12]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[26]) );
  DFFR_X1 constructing_unit_Datapath_diff_mult_h_int_samp_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_diff_mult_h_int[13]), .CK(clk), .RN(
        constructing_unit_Datapath_diff_mult_h_int_samp_n1), .Q(
        constructing_unit_Datapath_diff_mult_h_int[27]) );
  INV_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[0]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[11]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[1]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[12]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[2]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[13]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[3]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[14]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[4]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[15]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[5]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[16]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[6]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[17]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[7]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[18]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[8]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[19]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[9]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[20]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[21]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[22]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[23]) );
  DFFR_X1 constructing_unit_Datapath_MV0_int_v_ext_sample_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_MV0_int_v_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV0_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[24]) );
  XOR2_X1 constructing_unit_Datapath_R_sum_add_19_U2 ( .A(
        constructing_unit_Datapath_diff_mult_h_int[14]), .B(
        constructing_unit_Datapath_MV0_int_v_ext[11]), .Z(
        constructing_unit_Datapath_MV2p_int_v[0]) );
  AND2_X1 constructing_unit_Datapath_R_sum_add_19_U1 ( .A1(
        constructing_unit_Datapath_diff_mult_h_int[14]), .A2(
        constructing_unit_Datapath_MV0_int_v_ext[11]), .ZN(
        constructing_unit_Datapath_R_sum_add_19_n1) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_1 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[12]), .B(
        constructing_unit_Datapath_diff_mult_h_int[15]), .CI(
        constructing_unit_Datapath_R_sum_add_19_n1), .CO(
        constructing_unit_Datapath_R_sum_add_19_carry[2]), .S(
        constructing_unit_Datapath_MV2p_int_v[1]) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_2 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[13]), .B(
        constructing_unit_Datapath_diff_mult_h_int[16]), .CI(
        constructing_unit_Datapath_R_sum_add_19_carry[2]), .CO(
        constructing_unit_Datapath_R_sum_add_19_carry[3]), .S(
        constructing_unit_Datapath_MV2p_int_v[2]) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_3 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[14]), .B(
        constructing_unit_Datapath_diff_mult_h_int[17]), .CI(
        constructing_unit_Datapath_R_sum_add_19_carry[3]), .CO(
        constructing_unit_Datapath_R_sum_add_19_carry[4]), .S(
        constructing_unit_Datapath_MV2p_int_v[3]) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_4 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[15]), .B(
        constructing_unit_Datapath_diff_mult_h_int[18]), .CI(
        constructing_unit_Datapath_R_sum_add_19_carry[4]), .CO(
        constructing_unit_Datapath_R_sum_add_19_carry[5]), .S(
        constructing_unit_Datapath_MV2p_int_v[4]) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_5 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[16]), .B(
        constructing_unit_Datapath_diff_mult_h_int[19]), .CI(
        constructing_unit_Datapath_R_sum_add_19_carry[5]), .CO(
        constructing_unit_Datapath_R_sum_add_19_carry[6]), .S(
        constructing_unit_Datapath_MV2p_int_v[5]) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_6 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[17]), .B(
        constructing_unit_Datapath_diff_mult_h_int[20]), .CI(
        constructing_unit_Datapath_R_sum_add_19_carry[6]), .CO(
        constructing_unit_Datapath_R_sum_add_19_carry[7]), .S(
        constructing_unit_Datapath_MV2p_int_v[6]) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_7 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[18]), .B(
        constructing_unit_Datapath_diff_mult_h_int[21]), .CI(
        constructing_unit_Datapath_R_sum_add_19_carry[7]), .CO(
        constructing_unit_Datapath_R_sum_add_19_carry[8]), .S(
        constructing_unit_Datapath_MV2p_int_v[7]) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_8 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[19]), .B(
        constructing_unit_Datapath_diff_mult_h_int[22]), .CI(
        constructing_unit_Datapath_R_sum_add_19_carry[8]), .CO(
        constructing_unit_Datapath_R_sum_add_19_carry[9]), .S(
        constructing_unit_Datapath_MV2p_int_v[8]) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_9 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[20]), .B(
        constructing_unit_Datapath_diff_mult_h_int[23]), .CI(
        constructing_unit_Datapath_R_sum_add_19_carry[9]), .CO(
        constructing_unit_Datapath_R_sum_add_19_carry[10]), .S(
        constructing_unit_Datapath_MV2p_int_v[9]) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_10 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[21]), .B(
        constructing_unit_Datapath_diff_mult_h_int[24]), .CI(
        constructing_unit_Datapath_R_sum_add_19_carry[10]), .CO(
        constructing_unit_Datapath_R_sum_add_19_carry[11]), .S(
        constructing_unit_Datapath_MV2p_int_v[10]) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_11 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[22]), .B(
        constructing_unit_Datapath_diff_mult_h_int[25]), .CI(
        constructing_unit_Datapath_R_sum_add_19_carry[11]), .CO(
        constructing_unit_Datapath_R_sum_add_19_carry[12]), .S(
        constructing_unit_Datapath_MV2p_int_v[11]) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_12 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[23]), .B(
        constructing_unit_Datapath_diff_mult_h_int[26]), .CI(
        constructing_unit_Datapath_R_sum_add_19_carry[12]), .CO(
        constructing_unit_Datapath_R_sum_add_19_carry[13]), .S(
        constructing_unit_Datapath_MV2p_int_v[12]) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_13 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[24]), .B(
        constructing_unit_Datapath_diff_mult_h_int[27]), .CI(
        constructing_unit_Datapath_R_sum_add_19_carry[13]), .CO(
        constructing_unit_Datapath_R_sum_add_19_carry[14]), .S(
        constructing_unit_Datapath_MV2p_int_v[13]) );
  FA_X1 constructing_unit_Datapath_R_sum_add_19_U1_14 ( .A(
        constructing_unit_Datapath_MV0_int_v_ext[24]), .B(
        constructing_unit_Datapath_diff_mult_h_int[27]), .CI(
        constructing_unit_Datapath_R_sum_add_19_carry[14]), .S(
        constructing_unit_Datapath_MV2p_int_v[14]) );
  INV_X1 constructing_unit_Datapath_MV2p_int_v_sample_U4 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_MV2p_int_v_sample_n2) );
  INV_X1 constructing_unit_Datapath_MV2p_int_v_sample_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_MV2p_int_v_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[0]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_v[15]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[1]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_v[16]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[2]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_v[17]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[3]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_v[18]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[4]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_v[19]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[5]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_v[20]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[6]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_v[21]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[7]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_v[22]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[8]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_v[23]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[9]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_v[24]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_v[25]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[11]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n1), .Q(
        constructing_unit_Datapath_MV2p_int_v[26]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[12]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n2), .Q(
        constructing_unit_Datapath_MV2p_int_v[27]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[13]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n2), .Q(
        constructing_unit_Datapath_MV2p_int_v[28]) );
  DFFR_X1 constructing_unit_Datapath_MV2p_int_v_sample_Q_int_reg_14_ ( .D(
        constructing_unit_Datapath_MV2p_int_v[14]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2p_int_v_sample_n2), .Q(
        constructing_unit_Datapath_MV2p_int_v[29]) );
  INV_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_U4 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n2) );
  INV_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[0]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[11]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[1]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[12]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[2]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[13]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[3]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[14]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[4]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[15]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[5]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[16]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[6]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[17]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[7]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[18]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[8]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[19]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[9]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[20]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[21]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n1), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[22]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n2), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[23]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n2), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[24]) );
  DFFR_X1 constructing_unit_Datapath_MV2_int_v_ext_sample_Q_int_reg_14_ ( .D(
        constructing_unit_Datapath_MV2_int_v_ext[10]), .CK(clk), .RN(
        constructing_unit_Datapath_MV2_int_v_ext_sample_n2), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[25]) );
  XNOR2_X1 constructing_unit_Datapath_R_subD_sub_19_U18 ( .A(
        constructing_unit_Datapath_R_subD_sub_19_n16), .B(
        constructing_unit_Datapath_MV2p_int_v[15]), .ZN(
        constructing_unit_Datapath_D_v_tmp[0]) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U17 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[11]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n16) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U16 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[25]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n2) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U15 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[24]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n3) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U14 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[23]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n4) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U13 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[22]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n5) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U12 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[21]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n6) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U11 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[20]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n7) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U10 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[19]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n8) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U9 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[18]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n9) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U8 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[17]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n10) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U7 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[16]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n11) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U6 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[15]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n12) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U5 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[14]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n13) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U4 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[13]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n14) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U3 ( .A(
        constructing_unit_Datapath_MV2p_int_v[15]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n1) );
  NAND2_X1 constructing_unit_Datapath_R_subD_sub_19_U2 ( .A1(
        constructing_unit_Datapath_MV2_int_v_ext[11]), .A2(
        constructing_unit_Datapath_R_subD_sub_19_n1), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_carry[1]) );
  INV_X1 constructing_unit_Datapath_R_subD_sub_19_U1 ( .A(
        constructing_unit_Datapath_MV2_int_v_ext[12]), .ZN(
        constructing_unit_Datapath_R_subD_sub_19_n15) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_1 ( .A(
        constructing_unit_Datapath_MV2p_int_v[16]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n15), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[1]), .CO(
        constructing_unit_Datapath_R_subD_sub_19_carry[2]), .S(
        constructing_unit_Datapath_D_v_tmp[1]) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_2 ( .A(
        constructing_unit_Datapath_MV2p_int_v[17]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n14), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[2]), .CO(
        constructing_unit_Datapath_R_subD_sub_19_carry[3]), .S(
        constructing_unit_Datapath_D_v_tmp[2]) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_3 ( .A(
        constructing_unit_Datapath_MV2p_int_v[18]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n13), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[3]), .CO(
        constructing_unit_Datapath_R_subD_sub_19_carry[4]), .S(
        constructing_unit_Datapath_D_v_tmp[3]) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_4 ( .A(
        constructing_unit_Datapath_MV2p_int_v[19]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n12), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[4]), .CO(
        constructing_unit_Datapath_R_subD_sub_19_carry[5]), .S(
        constructing_unit_Datapath_D_v_tmp[4]) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_5 ( .A(
        constructing_unit_Datapath_MV2p_int_v[20]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n11), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[5]), .CO(
        constructing_unit_Datapath_R_subD_sub_19_carry[6]), .S(
        constructing_unit_Datapath_D_v_tmp[5]) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_6 ( .A(
        constructing_unit_Datapath_MV2p_int_v[21]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n10), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[6]), .CO(
        constructing_unit_Datapath_R_subD_sub_19_carry[7]), .S(
        constructing_unit_Datapath_D_v_tmp[6]) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_7 ( .A(
        constructing_unit_Datapath_MV2p_int_v[22]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n9), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[7]), .CO(
        constructing_unit_Datapath_R_subD_sub_19_carry[8]), .S(
        constructing_unit_Datapath_D_v_tmp[7]) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_8 ( .A(
        constructing_unit_Datapath_MV2p_int_v[23]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n8), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[8]), .CO(
        constructing_unit_Datapath_R_subD_sub_19_carry[9]), .S(
        constructing_unit_Datapath_D_v_tmp[8]) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_9 ( .A(
        constructing_unit_Datapath_MV2p_int_v[24]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n7), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[9]), .CO(
        constructing_unit_Datapath_R_subD_sub_19_carry[10]), .S(
        constructing_unit_Datapath_D_v_tmp[9]) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_10 ( .A(
        constructing_unit_Datapath_MV2p_int_v[25]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n6), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[10]), .CO(
        constructing_unit_Datapath_R_subD_sub_19_carry[11]), .S(
        constructing_unit_Datapath_D_v_tmp[10]) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_11 ( .A(
        constructing_unit_Datapath_MV2p_int_v[26]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n5), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[11]), .CO(
        constructing_unit_Datapath_R_subD_sub_19_carry[12]), .S(
        constructing_unit_Datapath_D_v_tmp[11]) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_12 ( .A(
        constructing_unit_Datapath_MV2p_int_v[27]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n4), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[12]), .CO(
        constructing_unit_Datapath_R_subD_sub_19_carry[13]), .S(
        constructing_unit_Datapath_D_v_tmp[12]) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_13 ( .A(
        constructing_unit_Datapath_MV2p_int_v[28]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n3), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[13]), .CO(
        constructing_unit_Datapath_R_subD_sub_19_carry[14]), .S(
        constructing_unit_Datapath_D_v_tmp[13]) );
  FA_X1 constructing_unit_Datapath_R_subD_sub_19_U2_14 ( .A(
        constructing_unit_Datapath_MV2p_int_v[29]), .B(
        constructing_unit_Datapath_R_subD_sub_19_n2), .CI(
        constructing_unit_Datapath_R_subD_sub_19_carry[14]), .S(
        constructing_unit_Datapath_D_v_tmp[14]) );
  INV_X1 constructing_unit_Datapath_D_v_sample_U4 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_D_v_sample_n2) );
  INV_X1 constructing_unit_Datapath_D_v_sample_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_D_v_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_D_v_tmp[0]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n1), .Q(
        constructing_unit_Datapath_D_v_0_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_D_v_tmp[1]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n1), .Q(
        constructing_unit_Datapath_D_v_1_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_D_v_tmp[2]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n1), .Q(
        constructing_unit_Datapath_D_v_2_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_D_v_tmp[3]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n1), .Q(
        constructing_unit_Datapath_D_v_3_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_D_v_tmp[4]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n1), .Q(
        constructing_unit_Datapath_D_v_4_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_D_v_tmp[5]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n1), .Q(
        constructing_unit_Datapath_D_v_5_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_D_v_tmp[6]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n1), .Q(
        constructing_unit_Datapath_D_v_6_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_D_v_tmp[7]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n1), .Q(
        constructing_unit_Datapath_D_v_7_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_D_v_tmp[8]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n1), .Q(
        constructing_unit_Datapath_D_v_8_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_D_v_tmp[9]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n1), .Q(
        constructing_unit_Datapath_D_v_9_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_D_v_tmp[10]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n1), .Q(
        constructing_unit_Datapath_D_v_10_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_D_v_tmp[11]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n1), .Q(
        constructing_unit_Datapath_D_v_11_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_D_v_tmp[12]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n2), .Q(
        constructing_unit_Datapath_D_v_12_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_D_v_tmp[13]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n2), .Q(
        constructing_unit_Datapath_D_v_13_) );
  DFFR_X1 constructing_unit_Datapath_D_v_sample_Q_int_reg_14_ ( .D(
        constructing_unit_Datapath_D_v_tmp[14]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sample_n2), .Q(
        constructing_unit_Datapath_D_v_14_) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U826 ( .A(
        constructing_unit_Datapath_D_v_13_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n776) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U825 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n666), .B(
        constructing_unit_Datapath_D_v_6_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n848) );
  NAND2_X1 constructing_unit_Datapath_R_squarer_mult_13_U824 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n848), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n763) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U823 ( .A(
        constructing_unit_Datapath_n16), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n778) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U822 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n776), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n778), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n112) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U821 ( .A(
        constructing_unit_Datapath_D_v_13_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n758) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U820 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n664), .B(
        constructing_unit_Datapath_D_v_4_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n847) );
  NAND2_X1 constructing_unit_Datapath_R_squarer_mult_13_U819 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n847), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n745) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U818 ( .A(
        constructing_unit_Datapath_n16), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n760) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U817 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n758), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n760), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n134) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U816 ( .A(
        constructing_unit_Datapath_D_v_13_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n740) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U815 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n662), .B(
        constructing_unit_Datapath_D_v_2_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n846) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U814 ( .A(
        constructing_unit_Datapath_n16), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n742) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U813 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n740), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n742), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n160) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U812 ( .A(
        constructing_unit_Datapath_D_v_2_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n809) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U811 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n672), .B(
        constructing_unit_Datapath_D_v_12_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n845) );
  NAND2_X1 constructing_unit_Datapath_R_squarer_mult_13_U810 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n845), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n706) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U809 ( .A(
        constructing_unit_Datapath_D_v_3_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n810) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U808 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n809), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n810), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n844) );
  XOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U807 ( .A(
        constructing_unit_Datapath_D_v_1_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n674), .Z(
        constructing_unit_Datapath_R_squarer_mult_13_n843) );
  NAND2_X1 constructing_unit_Datapath_R_squarer_mult_13_U806 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n843), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n689), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n842) );
  NAND2_X1 constructing_unit_Datapath_R_squarer_mult_13_U805 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n690), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n842), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n174) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U804 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n842), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n690), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n175) );
  AND3_X1 constructing_unit_Datapath_R_squarer_mult_13_U803 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n674), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n691), .A3(
        constructing_unit_Datapath_R_squarer_mult_13_n689), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n284) );
  OR3_X1 constructing_unit_Datapath_R_squarer_mult_13_U802 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .A2(
        constructing_unit_Datapath_D_v_0_), .A3(
        constructing_unit_Datapath_R_squarer_mult_13_n672), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n841) );
  OAI21_X1 constructing_unit_Datapath_R_squarer_mult_13_U801 ( .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n672), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .A(
        constructing_unit_Datapath_R_squarer_mult_13_n841), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n285) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U800 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n670), .B(
        constructing_unit_Datapath_D_v_10_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n840) );
  NAND2_X1 constructing_unit_Datapath_R_squarer_mult_13_U799 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n840), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n702) );
  OR3_X1 constructing_unit_Datapath_R_squarer_mult_13_U798 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .A2(
        constructing_unit_Datapath_D_v_0_), .A3(
        constructing_unit_Datapath_R_squarer_mult_13_n670), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n839) );
  OAI21_X1 constructing_unit_Datapath_R_squarer_mult_13_U797 ( .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n670), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .A(
        constructing_unit_Datapath_R_squarer_mult_13_n839), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n286) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U796 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n668), .B(
        constructing_unit_Datapath_D_v_8_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n838) );
  NAND2_X1 constructing_unit_Datapath_R_squarer_mult_13_U795 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n838), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n698) );
  OR3_X1 constructing_unit_Datapath_R_squarer_mult_13_U794 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .A2(
        constructing_unit_Datapath_D_v_0_), .A3(
        constructing_unit_Datapath_R_squarer_mult_13_n668), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n837) );
  OAI21_X1 constructing_unit_Datapath_R_squarer_mult_13_U793 ( .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n668), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .A(
        constructing_unit_Datapath_R_squarer_mult_13_n837), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n287) );
  OR3_X1 constructing_unit_Datapath_R_squarer_mult_13_U792 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .A2(
        constructing_unit_Datapath_D_v_0_), .A3(
        constructing_unit_Datapath_R_squarer_mult_13_n666), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n836) );
  OAI21_X1 constructing_unit_Datapath_R_squarer_mult_13_U791 ( .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n666), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .A(
        constructing_unit_Datapath_R_squarer_mult_13_n836), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n288) );
  OR3_X1 constructing_unit_Datapath_R_squarer_mult_13_U790 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .A2(
        constructing_unit_Datapath_D_v_0_), .A3(
        constructing_unit_Datapath_R_squarer_mult_13_n664), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n835) );
  OAI21_X1 constructing_unit_Datapath_R_squarer_mult_13_U789 ( .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n664), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .A(
        constructing_unit_Datapath_R_squarer_mult_13_n835), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n289) );
  OR3_X1 constructing_unit_Datapath_R_squarer_mult_13_U788 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .A2(
        constructing_unit_Datapath_D_v_0_), .A3(
        constructing_unit_Datapath_R_squarer_mult_13_n662), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n834) );
  OAI21_X1 constructing_unit_Datapath_R_squarer_mult_13_U787 ( .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n662), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .A(
        constructing_unit_Datapath_R_squarer_mult_13_n834), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n290) );
  NAND2_X1 constructing_unit_Datapath_R_squarer_mult_13_U786 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n709) );
  OAI21_X1 constructing_unit_Datapath_R_squarer_mult_13_U785 ( .B1(
        constructing_unit_Datapath_D_v_0_), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n660), .A(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n291) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U784 ( .A(
        constructing_unit_Datapath_D_v_13_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n833) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U783 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n833), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n293) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U782 ( .A(
        constructing_unit_Datapath_D_v_12_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n832) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U781 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n832), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n294) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U780 ( .A(
        constructing_unit_Datapath_D_v_11_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n831) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U779 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n831), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n295) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U778 ( .A(
        constructing_unit_Datapath_D_v_10_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n830) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U777 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n830), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n296) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U776 ( .A(
        constructing_unit_Datapath_D_v_9_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n829) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U775 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n829), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n297) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U774 ( .A(
        constructing_unit_Datapath_D_v_8_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n828) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U773 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n828), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n298) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U772 ( .A(
        constructing_unit_Datapath_D_v_7_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n827) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U771 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n827), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n299) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U770 ( .A(
        constructing_unit_Datapath_D_v_6_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n826) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U769 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n826), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n300) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U768 ( .A(
        constructing_unit_Datapath_D_v_5_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n825) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U767 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n825), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n301) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U766 ( .A(
        constructing_unit_Datapath_D_v_4_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n824) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U765 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n824), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n302) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U764 ( .A(
        constructing_unit_Datapath_D_v_3_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n823) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U763 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n823), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n303) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U762 ( .A(
        constructing_unit_Datapath_D_v_2_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n673), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n822) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U761 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n822), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n304) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U760 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n691), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n306) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U759 ( .A(
        constructing_unit_Datapath_n16), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n708) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U758 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n708), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n708), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n820) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U757 ( .A(
        constructing_unit_Datapath_D_v_12_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n819) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U756 ( .A(
        constructing_unit_Datapath_D_v_13_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n705) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U755 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n819), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n705), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n308) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U754 ( .A(
        constructing_unit_Datapath_D_v_11_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n818) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U753 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n818), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n819), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n309) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U752 ( .A(
        constructing_unit_Datapath_D_v_10_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n817) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U751 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n817), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n818), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n310) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U750 ( .A(
        constructing_unit_Datapath_D_v_9_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n816) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U749 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n816), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n817), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n311) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U748 ( .A(
        constructing_unit_Datapath_D_v_8_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n815) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U747 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n815), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n816), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n312) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U746 ( .A(
        constructing_unit_Datapath_D_v_7_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n814) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U745 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n814), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n815), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n313) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U744 ( .A(
        constructing_unit_Datapath_D_v_6_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n813) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U743 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n813), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n814), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n314) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U742 ( .A(
        constructing_unit_Datapath_D_v_5_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n812) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U741 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n812), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n813), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n315) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U740 ( .A(
        constructing_unit_Datapath_D_v_4_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n811) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U739 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n811), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n812), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n316) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U738 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n810), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n811), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n317) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U737 ( .A(
        constructing_unit_Datapath_D_v_1_), .B(
        constructing_unit_Datapath_D_v_13_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n808) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U736 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n808), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n809), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n319) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U735 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n671), .B(
        constructing_unit_Datapath_D_v_0_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n807) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U734 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n807), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n808), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n320) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U733 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n691), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n321) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U732 ( .A(
        constructing_unit_Datapath_n16), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n704) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U731 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n704), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n704), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n806) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U730 ( .A(
        constructing_unit_Datapath_D_v_12_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n805) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U729 ( .A(
        constructing_unit_Datapath_D_v_13_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n701) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U728 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n805), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n701), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n323) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U727 ( .A(
        constructing_unit_Datapath_D_v_11_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n804) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U726 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n804), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n805), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n324) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U725 ( .A(
        constructing_unit_Datapath_D_v_10_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n803) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U724 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n803), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n804), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n325) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U723 ( .A(
        constructing_unit_Datapath_D_v_9_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n802) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U722 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n802), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n803), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n326) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U721 ( .A(
        constructing_unit_Datapath_D_v_8_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n801) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U720 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n801), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n802), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n327) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U719 ( .A(
        constructing_unit_Datapath_D_v_7_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n800) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U718 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n800), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n801), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n328) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U717 ( .A(
        constructing_unit_Datapath_D_v_6_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n799) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U716 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n799), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n800), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n329) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U715 ( .A(
        constructing_unit_Datapath_D_v_5_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n798) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U714 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n798), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n799), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n330) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U713 ( .A(
        constructing_unit_Datapath_D_v_4_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n797) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U712 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n797), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n798), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n331) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U711 ( .A(
        constructing_unit_Datapath_D_v_3_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n796) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U710 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n796), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n797), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n332) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U709 ( .A(
        constructing_unit_Datapath_D_v_2_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n795) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U708 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n795), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n796), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n333) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U707 ( .A(
        constructing_unit_Datapath_D_v_1_), .B(
        constructing_unit_Datapath_D_v_11_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n794) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U706 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n794), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n795), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n334) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U705 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n669), .B(
        constructing_unit_Datapath_D_v_0_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n793) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U704 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n793), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n794), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n335) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U703 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n691), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n336) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U702 ( .A(
        constructing_unit_Datapath_n16), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n700) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U701 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n700), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n700), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n792) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U700 ( .A(
        constructing_unit_Datapath_D_v_12_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n791) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U699 ( .A(
        constructing_unit_Datapath_D_v_13_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n697) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U698 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n791), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n697), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n338) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U697 ( .A(
        constructing_unit_Datapath_D_v_11_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n790) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U696 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n790), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n791), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n339) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U695 ( .A(
        constructing_unit_Datapath_D_v_10_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n789) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U694 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n789), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n790), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n340) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U693 ( .A(
        constructing_unit_Datapath_D_v_9_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n788) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U692 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n788), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n789), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n341) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U691 ( .A(
        constructing_unit_Datapath_D_v_8_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n787) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U690 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n787), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n788), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n342) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U689 ( .A(
        constructing_unit_Datapath_D_v_7_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n786) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U688 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n786), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n787), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n343) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U687 ( .A(
        constructing_unit_Datapath_D_v_6_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n785) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U686 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n785), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n786), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n344) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U685 ( .A(
        constructing_unit_Datapath_D_v_5_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n784) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U684 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n784), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n785), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n345) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U683 ( .A(
        constructing_unit_Datapath_D_v_4_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n783) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U682 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n783), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n784), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n346) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U681 ( .A(
        constructing_unit_Datapath_D_v_3_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n782) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U680 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n782), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n783), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n347) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U679 ( .A(
        constructing_unit_Datapath_D_v_2_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n781) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U678 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n781), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n782), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n348) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U677 ( .A(
        constructing_unit_Datapath_D_v_1_), .B(
        constructing_unit_Datapath_D_v_9_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n780) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U676 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n780), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n781), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n349) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U675 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n667), .B(
        constructing_unit_Datapath_D_v_0_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n779) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U674 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n779), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n780), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n350) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U673 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n691), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n351) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U672 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n778), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n778), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n777) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U671 ( .A(
        constructing_unit_Datapath_D_v_12_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n775) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U670 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n775), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n776), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n353) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U669 ( .A(
        constructing_unit_Datapath_D_v_11_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n774) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U668 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n774), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n775), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n354) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U667 ( .A(
        constructing_unit_Datapath_D_v_10_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n773) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U666 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n773), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n774), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n355) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U665 ( .A(
        constructing_unit_Datapath_D_v_9_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n772) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U664 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n772), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n773), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n356) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U663 ( .A(
        constructing_unit_Datapath_D_v_8_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n771) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U662 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n771), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n772), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n357) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U661 ( .A(
        constructing_unit_Datapath_D_v_7_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n770) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U660 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n770), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n771), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n358) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U659 ( .A(
        constructing_unit_Datapath_D_v_6_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n769) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U658 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n769), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n770), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n359) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U657 ( .A(
        constructing_unit_Datapath_D_v_5_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n768) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U656 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n768), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n769), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n360) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U655 ( .A(
        constructing_unit_Datapath_D_v_4_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n767) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U654 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n767), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n768), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n361) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U653 ( .A(
        constructing_unit_Datapath_D_v_3_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n766) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U652 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n766), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n767), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n362) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U651 ( .A(
        constructing_unit_Datapath_D_v_2_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n765) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U650 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n765), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n766), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n363) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U649 ( .A(
        constructing_unit_Datapath_D_v_1_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n764) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U648 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n764), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n765), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n364) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U647 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n665), .B(
        constructing_unit_Datapath_D_v_0_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n762) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U646 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n762), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n763), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n764), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n365) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U645 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n691), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n761), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n366) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U644 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n760), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n760), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n759) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U643 ( .A(
        constructing_unit_Datapath_D_v_12_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n757) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U642 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n757), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n758), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n368) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U641 ( .A(
        constructing_unit_Datapath_D_v_11_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n756) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U640 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n756), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n757), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n369) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U639 ( .A(
        constructing_unit_Datapath_D_v_10_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n755) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U638 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n755), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n756), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n370) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U637 ( .A(
        constructing_unit_Datapath_D_v_9_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n754) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U636 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n754), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n755), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n371) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U635 ( .A(
        constructing_unit_Datapath_D_v_8_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n753) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U634 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n753), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n754), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n372) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U633 ( .A(
        constructing_unit_Datapath_D_v_7_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n752) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U632 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n752), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n753), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n373) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U631 ( .A(
        constructing_unit_Datapath_D_v_6_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n751) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U630 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n751), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n752), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n374) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U629 ( .A(
        constructing_unit_Datapath_D_v_5_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n750) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U628 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n750), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n751), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n375) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U627 ( .A(
        constructing_unit_Datapath_D_v_4_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n749) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U626 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n749), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n750), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n376) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U625 ( .A(
        constructing_unit_Datapath_D_v_3_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n748) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U624 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n748), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n749), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n377) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U623 ( .A(
        constructing_unit_Datapath_D_v_2_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n747) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U622 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n747), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n748), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n378) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U621 ( .A(
        constructing_unit_Datapath_D_v_1_), .B(
        constructing_unit_Datapath_D_v_5_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n746) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U620 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n746), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n747), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n379) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U619 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n663), .B(
        constructing_unit_Datapath_D_v_0_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n744) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U618 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n744), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n745), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n746), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n380) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U617 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n691), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n743), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n381) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U616 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n742), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n742), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n741) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U615 ( .A(
        constructing_unit_Datapath_D_v_12_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n739) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U614 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n739), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n740), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n383) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U613 ( .A(
        constructing_unit_Datapath_D_v_11_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n738) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U612 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n738), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n739), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n384) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U611 ( .A(
        constructing_unit_Datapath_D_v_10_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n737) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U610 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n737), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n738), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n385) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U609 ( .A(
        constructing_unit_Datapath_D_v_9_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n736) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U608 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n736), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n737), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n386) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U607 ( .A(
        constructing_unit_Datapath_D_v_8_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n735) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U606 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n735), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n736), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n387) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U605 ( .A(
        constructing_unit_Datapath_D_v_7_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n734) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U604 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n734), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n735), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n388) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U603 ( .A(
        constructing_unit_Datapath_D_v_6_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n733) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U602 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n733), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n734), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n389) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U601 ( .A(
        constructing_unit_Datapath_D_v_5_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n732) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U600 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n732), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n733), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n390) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U599 ( .A(
        constructing_unit_Datapath_D_v_4_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n731) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U598 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n731), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n732), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n391) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U597 ( .A(
        constructing_unit_Datapath_D_v_3_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n730) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U596 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n730), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n731), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n392) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U595 ( .A(
        constructing_unit_Datapath_D_v_2_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n729) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U594 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n729), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n730), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n393) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U593 ( .A(
        constructing_unit_Datapath_D_v_1_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n728) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U592 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n728), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n729), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n394) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U591 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n661), .B(
        constructing_unit_Datapath_D_v_0_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n726) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U590 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n726), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n727), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n728), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n395) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U589 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n691), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n396) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U588 ( .A(
        constructing_unit_Datapath_n16), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n723) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U587 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n723), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n723), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n724) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U586 ( .A(
        constructing_unit_Datapath_D_v_13_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n722) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U585 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n722), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n723), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n398) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U584 ( .A(
        constructing_unit_Datapath_D_v_12_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n721) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U583 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n721), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n722), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n399) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U582 ( .A(
        constructing_unit_Datapath_D_v_11_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n720) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U581 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n720), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n721), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n400) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U580 ( .A(
        constructing_unit_Datapath_D_v_10_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n719) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U579 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n719), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n720), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n401) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U578 ( .A(
        constructing_unit_Datapath_D_v_9_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n718) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U577 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n718), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n719), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n402) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U576 ( .A(
        constructing_unit_Datapath_D_v_8_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n717) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U575 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n717), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n718), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n403) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U574 ( .A(
        constructing_unit_Datapath_D_v_7_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n716) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U573 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n716), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n717), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n404) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U572 ( .A(
        constructing_unit_Datapath_D_v_6_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n715) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U571 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n715), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n716), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n405) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U570 ( .A(
        constructing_unit_Datapath_D_v_5_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n714) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U569 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n714), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n715), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n406) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U568 ( .A(
        constructing_unit_Datapath_D_v_4_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n713) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U567 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n713), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n714), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n407) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U566 ( .A(
        constructing_unit_Datapath_D_v_3_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n712) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U565 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n712), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n713), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n408) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U564 ( .A(
        constructing_unit_Datapath_D_v_2_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n711) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U563 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n711), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n712), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n409) );
  XNOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U562 ( .A(
        constructing_unit_Datapath_D_v_1_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n659), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n710) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U561 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n710), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n711), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n410) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U560 ( .A1(
        constructing_unit_Datapath_D_v_0_), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n709), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n710), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n411) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U559 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n705), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n706), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n707), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n708), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n70) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U558 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n701), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n702), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n703), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n704), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n80) );
  OAI22_X1 constructing_unit_Datapath_R_squarer_mult_13_U557 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n697), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n698), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n699), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n700), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n94) );
  NOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U556 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n691), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n692), .ZN(
        constructing_unit_Datapath_D_v_sq_tmp[0]) );
  XOR2_X1 constructing_unit_Datapath_R_squarer_mult_13_U555 ( .A(
        constructing_unit_Datapath_n16), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n674), .Z(
        constructing_unit_Datapath_R_squarer_mult_13_n696) );
  NAND2_X1 constructing_unit_Datapath_R_squarer_mult_13_U554 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n696), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n689), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n693) );
  AOI222_X1 constructing_unit_Datapath_R_squarer_mult_13_U553 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n38), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n68), .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n38), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n67), .C1(
        constructing_unit_Datapath_R_squarer_mult_13_n67), .C2(
        constructing_unit_Datapath_R_squarer_mult_13_n68), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n695) );
  AND2_X1 constructing_unit_Datapath_R_squarer_mult_13_U552 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n693), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n675), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n694) );
  AOI221_X1 constructing_unit_Datapath_R_squarer_mult_13_U551 ( .B1(
        constructing_unit_Datapath_R_squarer_mult_13_n66), .B2(
        constructing_unit_Datapath_R_squarer_mult_13_n693), .C1(
        constructing_unit_Datapath_R_squarer_mult_13_n66), .C2(
        constructing_unit_Datapath_R_squarer_mult_13_n675), .A(
        constructing_unit_Datapath_R_squarer_mult_13_n694), .ZN(
        constructing_unit_Datapath_R_squarer_product_29_) );
  INV_X2 constructing_unit_Datapath_R_squarer_mult_13_U550 ( .A(
        constructing_unit_Datapath_D_v_0_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n692) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U549 ( .A(
        constructing_unit_Datapath_D_v_13_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n672) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U548 ( .A(
        constructing_unit_Datapath_D_v_11_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n670) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U547 ( .A(
        constructing_unit_Datapath_D_v_9_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n668) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U546 ( .A(
        constructing_unit_Datapath_D_v_7_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n666) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U545 ( .A(
        constructing_unit_Datapath_D_v_5_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n664) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U544 ( .A(
        constructing_unit_Datapath_D_v_3_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n662) );
  XOR2_X2 constructing_unit_Datapath_R_squarer_mult_13_U543 ( .A(
        constructing_unit_Datapath_D_v_6_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n664), .Z(
        constructing_unit_Datapath_R_squarer_mult_13_n761) );
  XOR2_X2 constructing_unit_Datapath_R_squarer_mult_13_U542 ( .A(
        constructing_unit_Datapath_D_v_4_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n662), .Z(
        constructing_unit_Datapath_R_squarer_mult_13_n743) );
  XOR2_X2 constructing_unit_Datapath_R_squarer_mult_13_U541 ( .A(
        constructing_unit_Datapath_D_v_2_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n660), .Z(
        constructing_unit_Datapath_R_squarer_mult_13_n725) );
  XOR2_X2 constructing_unit_Datapath_R_squarer_mult_13_U540 ( .A(
        constructing_unit_Datapath_D_v_12_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n670), .Z(
        constructing_unit_Datapath_R_squarer_mult_13_n707) );
  XOR2_X2 constructing_unit_Datapath_R_squarer_mult_13_U539 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n674), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n672), .Z(
        constructing_unit_Datapath_R_squarer_mult_13_n821) );
  XOR2_X2 constructing_unit_Datapath_R_squarer_mult_13_U538 ( .A(
        constructing_unit_Datapath_D_v_10_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n668), .Z(
        constructing_unit_Datapath_R_squarer_mult_13_n703) );
  XOR2_X2 constructing_unit_Datapath_R_squarer_mult_13_U537 ( .A(
        constructing_unit_Datapath_D_v_8_), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n666), .Z(
        constructing_unit_Datapath_R_squarer_mult_13_n699) );
  INV_X2 constructing_unit_Datapath_R_squarer_mult_13_U536 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n660), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n659) );
  NAND2_X2 constructing_unit_Datapath_R_squarer_mult_13_U535 ( .A1(
        constructing_unit_Datapath_R_squarer_mult_13_n725), .A2(
        constructing_unit_Datapath_R_squarer_mult_13_n846), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n727) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U534 ( .A(
        constructing_unit_Datapath_D_v_1_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n660) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U533 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n70), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n682) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U532 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n759), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n686) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U531 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n741), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n684) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U530 ( .A(
        constructing_unit_Datapath_D_v_0_), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n691) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U529 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n695), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n675) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U528 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n820), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n681) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U527 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n806), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n679) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U526 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n777), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n688) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U525 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n112), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n687) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U524 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n792), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n677) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U523 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n80), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n680) );
  BUF_X1 constructing_unit_Datapath_R_squarer_mult_13_U522 ( .A(
        constructing_unit_Datapath_n16), .Z(
        constructing_unit_Datapath_R_squarer_mult_13_n673) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U521 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n844), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n690) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U520 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n134), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n685) );
  BUF_X1 constructing_unit_Datapath_R_squarer_mult_13_U519 ( .A(
        constructing_unit_Datapath_n16), .Z(
        constructing_unit_Datapath_R_squarer_mult_13_n674) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U518 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n160), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n683) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U517 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n724), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n676) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U516 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n662), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n661) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U515 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n666), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n665) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U514 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n664), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n663) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U513 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n668), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n667) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U512 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n672), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n671) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U511 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n670), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n669) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U510 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n94), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n678) );
  INV_X1 constructing_unit_Datapath_R_squarer_mult_13_U509 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n821), .ZN(
        constructing_unit_Datapath_R_squarer_mult_13_n689) );
  HA_X1 constructing_unit_Datapath_R_squarer_mult_13_U163 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n395), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n409), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n258), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n259) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U162 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n408), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n381), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n394), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n256), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n257) );
  HA_X1 constructing_unit_Datapath_R_squarer_mult_13_U161 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n289), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n380), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n254), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n255) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U160 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n393), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n407), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n255), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n252), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n253) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U159 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n406), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n366), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n392), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n250), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n251) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U158 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n254), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n379), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n251), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n248), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n249) );
  HA_X1 constructing_unit_Datapath_R_squarer_mult_13_U157 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n288), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n365), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n246), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n247) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U156 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n378), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n405), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n391), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n244), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n245) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U155 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n250), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n247), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n245), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n242), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n243) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U154 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n377), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n351), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n404), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n240), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n241) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U153 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n364), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n390), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n246), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n238), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n239) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U152 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n241), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n244), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n239), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n236), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n237) );
  HA_X1 constructing_unit_Datapath_R_squarer_mult_13_U151 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n287), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n350), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n234), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n235) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U150 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n363), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n376), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n389), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n232), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n233) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U149 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n235), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n403), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n240), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n230), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n231) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U148 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n233), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n238), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n231), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n228), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n229) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U147 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n362), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n336), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n402), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n226), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n227) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U146 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n349), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n388), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n375), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n224), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n225) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U145 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n232), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n234), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n227), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n222), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n223) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U144 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n230), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n225), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n223), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n220), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n221) );
  HA_X1 constructing_unit_Datapath_R_squarer_mult_13_U143 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n286), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n335), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n218), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n219) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U142 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n348), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n374), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n401), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n216), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n217) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U141 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n361), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n387), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n219), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n214), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n215) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U140 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n224), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n226), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n217), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n212), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n213) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U139 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n222), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n215), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n213), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n210), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n211) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U138 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n347), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n321), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n400), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n208), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n209) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U137 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n334), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n386), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n360), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n206), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n207) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U136 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n218), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n373), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n216), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n204), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n205) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U135 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n207), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n209), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n214), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n202), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n203) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U134 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n205), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n212), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n203), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n200), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n201) );
  HA_X1 constructing_unit_Datapath_R_squarer_mult_13_U133 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n285), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n320), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n198), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n199) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U132 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n399), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n359), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n385), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n196), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n197) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U131 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n333), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n372), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n346), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n194), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n195) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U130 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n208), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n199), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n206), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n192), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n193) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U129 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n197), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n195), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n204), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n190), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n191) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U128 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n202), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n193), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n191), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n188), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n189) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U127 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n332), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n306), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n398), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n186), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n187) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U126 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n319), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n384), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n345), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n184), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n185) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U125 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n358), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n371), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n198), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n182), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n183) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U124 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n194), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n196), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n187), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n180), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n181) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U123 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n183), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n185), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n192), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n178), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n179) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U122 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n181), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n190), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n179), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n176), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n177) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U119 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n284), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n357), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n676), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n172), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n173) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U118 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n383), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n331), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n344), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n170), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n171) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U117 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n175), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n370), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n186), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n168), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n169) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U116 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n182), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n184), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n171), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n166), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n167) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U115 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n180), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n173), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n169), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n164), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n165) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U114 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n167), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n178), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n165), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n162), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n163) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U112 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n369), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n330), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n304), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n158), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n159) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U111 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n317), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n356), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n343), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n156), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n157) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U110 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n174), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n683), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n172), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n154), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n155) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U109 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n157), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n170), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n159), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n152), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n153) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U108 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n166), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n168), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n155), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n150), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n151) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U107 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n164), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n153), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n151), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n148), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n149) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U106 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n160), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n303), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n684), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n146), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n147) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U105 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n316), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n368), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n355), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n144), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n145) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U104 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n329), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n342), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n158), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n142), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n143) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U103 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n145), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n156), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n147), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n140), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n141) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U102 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n143), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n154), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n152), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n138), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n139) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U101 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n150), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n141), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n139), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n136), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n137) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U99 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n354), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n328), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n341), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n132), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n133) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U98 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n302), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n315), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n685), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n130), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n131) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U97 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n144), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n146), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n133), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n128), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n129) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U96 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n142), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n131), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n140), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n126), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n127) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U95 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n138), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n129), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n127), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n124), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n125) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U94 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n134), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n301), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n686), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n122), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n123) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U93 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n314), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n353), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n327), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n120), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n121) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U92 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n132), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n340), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n130), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n118), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n119) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U91 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n123), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n121), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n128), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n116), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n117) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U90 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n126), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n119), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n117), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n114), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n115) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U88 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n339), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n313), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n300), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n110), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n111) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U87 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n687), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n326), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n122), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n108), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n109) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U86 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n111), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n120), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n118), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n106), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n107) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U85 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n116), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n109), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n107), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n104), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n105) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U84 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n338), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n299), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n688), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n102), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n103) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U83 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n312), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n112), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n325), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n100), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n101) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U82 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n101), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n110), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n103), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n98), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n99) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U81 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n106), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n108), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n99), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n96), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n97) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U79 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n298), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n311), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n324), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n92), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n93) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U78 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n102), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n678), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n100), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n90), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n91) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U77 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n91), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n93), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n98), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n88), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n89) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U76 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n310), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n297), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n677), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n86), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n87) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U75 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n94), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n323), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n92), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n84), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n85) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U74 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n90), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n87), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n85), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n82), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n83) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U72 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n296), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n309), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n680), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n78), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n79) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U71 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n79), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n86), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n84), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n76), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n77) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U70 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n308), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n80), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n679), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n74), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n75) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U69 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n78), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n295), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n75), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n72), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n73) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U67 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n682), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n294), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n74), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n68), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n69) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U66 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n293), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n70), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n681), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n66), .S(
        constructing_unit_Datapath_R_squarer_mult_13_n67) );
  HA_X1 constructing_unit_Datapath_R_squarer_mult_13_U64 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n411), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n291), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n63), .S(
        constructing_unit_Datapath_D_v_sq_tmp[1]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U63 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n410), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n396), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n63), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n62), .S(
        constructing_unit_Datapath_D_v_sq_tmp[2]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U62 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n259), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n290), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n62), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n61), .S(
        constructing_unit_Datapath_D_v_sq_tmp[3]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U61 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n257), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n258), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n61), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n60), .S(
        constructing_unit_Datapath_D_v_sq_tmp[4]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U60 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n253), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n256), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n60), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n59), .S(
        constructing_unit_Datapath_D_v_sq_tmp[5]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U59 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n249), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n252), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n59), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n58), .S(
        constructing_unit_Datapath_D_v_sq_tmp[6]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U58 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n243), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n248), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n58), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n57), .S(
        constructing_unit_Datapath_D_v_sq_tmp[7]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U57 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n237), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n242), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n57), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n56), .S(
        constructing_unit_Datapath_D_v_sq_tmp[8]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U56 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n229), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n236), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n56), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n55), .S(
        constructing_unit_Datapath_D_v_sq_tmp[9]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U55 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n221), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n228), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n55), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n54), .S(
        constructing_unit_Datapath_D_v_sq_tmp[10]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U54 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n211), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n220), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n54), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n53), .S(
        constructing_unit_Datapath_D_v_sq_tmp[11]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U53 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n201), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n210), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n53), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n52), .S(
        constructing_unit_Datapath_D_v_sq_tmp[12]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U52 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n189), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n200), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n52), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n51), .S(
        constructing_unit_Datapath_D_v_sq_tmp[13]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U51 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n177), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n188), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n51), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n50), .S(
        constructing_unit_Datapath_D_v_sq_tmp[14]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U50 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n163), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n176), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n50), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n49), .S(
        constructing_unit_Datapath_D_v_sq_tmp[15]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U49 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n149), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n162), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n49), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n48), .S(
        constructing_unit_Datapath_D_v_sq_tmp[16]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U48 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n137), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n148), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n48), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n47), .S(
        constructing_unit_Datapath_D_v_sq_tmp[17]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U47 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n125), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n136), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n47), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n46), .S(
        constructing_unit_Datapath_D_v_sq_tmp[18]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U46 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n115), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n124), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n46), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n45), .S(
        constructing_unit_Datapath_D_v_sq_tmp[19]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U45 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n105), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n114), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n45), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n44), .S(
        constructing_unit_Datapath_D_v_sq_tmp[20]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U44 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n97), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n104), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n44), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n43), .S(
        constructing_unit_Datapath_D_v_sq_tmp[21]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U43 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n89), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n96), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n43), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n42), .S(
        constructing_unit_Datapath_D_v_sq_tmp[22]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U42 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n83), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n88), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n42), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n41), .S(
        constructing_unit_Datapath_D_v_sq_tmp[23]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U41 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n77), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n82), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n41), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n40), .S(
        constructing_unit_Datapath_D_v_sq_tmp[24]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U40 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n73), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n76), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n40), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n39), .S(
        constructing_unit_Datapath_D_v_sq_tmp[25]) );
  FA_X1 constructing_unit_Datapath_R_squarer_mult_13_U39 ( .A(
        constructing_unit_Datapath_R_squarer_mult_13_n69), .B(
        constructing_unit_Datapath_R_squarer_mult_13_n72), .CI(
        constructing_unit_Datapath_R_squarer_mult_13_n39), .CO(
        constructing_unit_Datapath_R_squarer_mult_13_n38), .S(
        constructing_unit_Datapath_D_v_sq_tmp[26]) );
  OR3_X1 constructing_unit_Datapath_MV0_check_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__9_), .A2(
        constructing_unit_Datapath_MV0_int_v_1__8_), .A3(
        constructing_unit_Datapath_MV0_int_v_1__7_), .ZN(
        constructing_unit_Datapath_MV0_check_n10) );
  OR3_X1 constructing_unit_Datapath_MV0_check_U10 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__9_), .A2(
        constructing_unit_Datapath_MV0_int_h_1__8_), .A3(
        constructing_unit_Datapath_MV0_int_h_1__7_), .ZN(
        constructing_unit_Datapath_MV0_check_n7) );
  NOR4_X1 constructing_unit_Datapath_MV0_check_U9 ( .A1(
        constructing_unit_Datapath_MV0_check_n10), .A2(
        constructing_unit_Datapath_MV0_int_v_1__4_), .A3(
        constructing_unit_Datapath_MV0_int_v_1__6_), .A4(
        constructing_unit_Datapath_MV0_int_v_1__5_), .ZN(
        constructing_unit_Datapath_MV0_check_n9) );
  NOR3_X1 constructing_unit_Datapath_MV0_check_U8 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__1_), .A2(
        constructing_unit_Datapath_MV0_int_v_1__3_), .A3(
        constructing_unit_Datapath_MV0_int_v_1__2_), .ZN(
        constructing_unit_Datapath_MV0_check_n8) );
  INV_X1 constructing_unit_Datapath_MV0_check_U7 ( .A(
        constructing_unit_Datapath_MV0_int_v_1__0_), .ZN(
        constructing_unit_Datapath_MV0_check_n2) );
  NAND4_X1 constructing_unit_Datapath_MV0_check_U6 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__10_), .A2(
        constructing_unit_Datapath_MV0_check_n2), .A3(
        constructing_unit_Datapath_MV0_check_n8), .A4(
        constructing_unit_Datapath_MV0_check_n9), .ZN(
        constructing_unit_Datapath_MV0_check_n3) );
  NOR4_X1 constructing_unit_Datapath_MV0_check_U5 ( .A1(
        constructing_unit_Datapath_MV0_check_n7), .A2(
        constructing_unit_Datapath_MV0_int_h_1__4_), .A3(
        constructing_unit_Datapath_MV0_int_h_1__6_), .A4(
        constructing_unit_Datapath_MV0_int_h_1__5_), .ZN(
        constructing_unit_Datapath_MV0_check_n6) );
  NOR3_X1 constructing_unit_Datapath_MV0_check_U4 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__1_), .A2(
        constructing_unit_Datapath_MV0_int_h_1__3_), .A3(
        constructing_unit_Datapath_MV0_int_h_1__2_), .ZN(
        constructing_unit_Datapath_MV0_check_n5) );
  INV_X1 constructing_unit_Datapath_MV0_check_U3 ( .A(
        constructing_unit_Datapath_MV0_int_h_1__0_), .ZN(
        constructing_unit_Datapath_MV0_check_n1) );
  NAND4_X1 constructing_unit_Datapath_MV0_check_U2 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__10_), .A2(
        constructing_unit_Datapath_MV0_check_n1), .A3(
        constructing_unit_Datapath_MV0_check_n5), .A4(
        constructing_unit_Datapath_MV0_check_n6), .ZN(
        constructing_unit_Datapath_MV0_check_n4) );
  NAND2_X1 constructing_unit_Datapath_MV0_check_U1 ( .A1(
        constructing_unit_Datapath_MV0_check_n3), .A2(
        constructing_unit_Datapath_MV0_check_n4), .ZN(
        constructing_unit_Datapath_UA_flag[0]) );
  OR3_X1 constructing_unit_Datapath_MV1_check_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__9_), .A2(
        constructing_unit_Datapath_MV1_int_v_1__8_), .A3(
        constructing_unit_Datapath_MV1_int_v_1__7_), .ZN(
        constructing_unit_Datapath_MV1_check_n11) );
  OR3_X1 constructing_unit_Datapath_MV1_check_U10 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__9_), .A2(
        constructing_unit_Datapath_MV1_int_h_1__8_), .A3(
        constructing_unit_Datapath_MV1_int_h_1__7_), .ZN(
        constructing_unit_Datapath_MV1_check_n14) );
  NOR4_X1 constructing_unit_Datapath_MV1_check_U9 ( .A1(
        constructing_unit_Datapath_MV1_check_n11), .A2(
        constructing_unit_Datapath_MV1_int_v_1__4_), .A3(
        constructing_unit_Datapath_MV1_int_v_1__6_), .A4(
        constructing_unit_Datapath_MV1_int_v_1__5_), .ZN(
        constructing_unit_Datapath_MV1_check_n12) );
  INV_X1 constructing_unit_Datapath_MV1_check_U8 ( .A(
        constructing_unit_Datapath_MV1_int_v_1__0_), .ZN(
        constructing_unit_Datapath_MV1_check_n1) );
  NOR3_X1 constructing_unit_Datapath_MV1_check_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__1_), .A2(
        constructing_unit_Datapath_MV1_int_v_1__3_), .A3(
        constructing_unit_Datapath_MV1_int_v_1__2_), .ZN(
        constructing_unit_Datapath_MV1_check_n13) );
  NAND4_X1 constructing_unit_Datapath_MV1_check_U6 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__10_), .A2(
        constructing_unit_Datapath_MV1_check_n1), .A3(
        constructing_unit_Datapath_MV1_check_n13), .A4(
        constructing_unit_Datapath_MV1_check_n12), .ZN(
        constructing_unit_Datapath_MV1_check_n18) );
  NOR4_X1 constructing_unit_Datapath_MV1_check_U5 ( .A1(
        constructing_unit_Datapath_MV1_check_n14), .A2(
        constructing_unit_Datapath_MV1_int_h_1__4_), .A3(
        constructing_unit_Datapath_MV1_int_h_1__6_), .A4(
        constructing_unit_Datapath_MV1_int_h_1__5_), .ZN(
        constructing_unit_Datapath_MV1_check_n15) );
  INV_X1 constructing_unit_Datapath_MV1_check_U4 ( .A(
        constructing_unit_Datapath_MV1_int_h_1__0_), .ZN(
        constructing_unit_Datapath_MV1_check_n2) );
  NOR3_X1 constructing_unit_Datapath_MV1_check_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__1_), .A2(
        constructing_unit_Datapath_MV1_int_h_1__3_), .A3(
        constructing_unit_Datapath_MV1_int_h_1__2_), .ZN(
        constructing_unit_Datapath_MV1_check_n16) );
  NAND4_X1 constructing_unit_Datapath_MV1_check_U2 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__10_), .A2(
        constructing_unit_Datapath_MV1_check_n2), .A3(
        constructing_unit_Datapath_MV1_check_n16), .A4(
        constructing_unit_Datapath_MV1_check_n15), .ZN(
        constructing_unit_Datapath_MV1_check_n17) );
  NAND2_X1 constructing_unit_Datapath_MV1_check_U1 ( .A1(
        constructing_unit_Datapath_MV1_check_n18), .A2(
        constructing_unit_Datapath_MV1_check_n17), .ZN(
        constructing_unit_Datapath_UA_flag[1]) );
  OR3_X1 constructing_unit_Datapath_MV2_check_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__9_), .A2(
        constructing_unit_Datapath_MV2_int_v_1__8_), .A3(
        constructing_unit_Datapath_MV2_int_v_1__7_), .ZN(
        constructing_unit_Datapath_MV2_check_n11) );
  OR3_X1 constructing_unit_Datapath_MV2_check_U10 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__9_), .A2(
        constructing_unit_Datapath_MV2_int_h_1__8_), .A3(
        constructing_unit_Datapath_MV2_int_h_1__7_), .ZN(
        constructing_unit_Datapath_MV2_check_n14) );
  NOR4_X1 constructing_unit_Datapath_MV2_check_U9 ( .A1(
        constructing_unit_Datapath_MV2_check_n11), .A2(
        constructing_unit_Datapath_MV2_int_v_1__4_), .A3(
        constructing_unit_Datapath_MV2_int_v_1__6_), .A4(
        constructing_unit_Datapath_MV2_int_v_1__5_), .ZN(
        constructing_unit_Datapath_MV2_check_n12) );
  NOR3_X1 constructing_unit_Datapath_MV2_check_U8 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__1_), .A2(
        constructing_unit_Datapath_MV2_int_v_1__3_), .A3(
        constructing_unit_Datapath_MV2_int_v_1__2_), .ZN(
        constructing_unit_Datapath_MV2_check_n13) );
  INV_X1 constructing_unit_Datapath_MV2_check_U7 ( .A(
        constructing_unit_Datapath_MV2_int_v_1__0_), .ZN(
        constructing_unit_Datapath_MV2_check_n1) );
  NAND4_X1 constructing_unit_Datapath_MV2_check_U6 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__10_), .A2(
        constructing_unit_Datapath_MV2_check_n1), .A3(
        constructing_unit_Datapath_MV2_check_n13), .A4(
        constructing_unit_Datapath_MV2_check_n12), .ZN(
        constructing_unit_Datapath_MV2_check_n18) );
  NOR4_X1 constructing_unit_Datapath_MV2_check_U5 ( .A1(
        constructing_unit_Datapath_MV2_check_n14), .A2(
        constructing_unit_Datapath_MV2_int_h_1__4_), .A3(
        constructing_unit_Datapath_MV2_int_h_1__6_), .A4(
        constructing_unit_Datapath_MV2_int_h_1__5_), .ZN(
        constructing_unit_Datapath_MV2_check_n15) );
  NOR3_X1 constructing_unit_Datapath_MV2_check_U4 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__1_), .A2(
        constructing_unit_Datapath_MV2_int_h_1__3_), .A3(
        constructing_unit_Datapath_MV2_int_h_1__2_), .ZN(
        constructing_unit_Datapath_MV2_check_n16) );
  INV_X1 constructing_unit_Datapath_MV2_check_U3 ( .A(
        constructing_unit_Datapath_MV2_int_h_1__0_), .ZN(
        constructing_unit_Datapath_MV2_check_n2) );
  NAND4_X1 constructing_unit_Datapath_MV2_check_U2 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__10_), .A2(
        constructing_unit_Datapath_MV2_check_n2), .A3(
        constructing_unit_Datapath_MV2_check_n16), .A4(
        constructing_unit_Datapath_MV2_check_n15), .ZN(
        constructing_unit_Datapath_MV2_check_n17) );
  NAND2_X1 constructing_unit_Datapath_MV2_check_U1 ( .A1(
        constructing_unit_Datapath_MV2_check_n18), .A2(
        constructing_unit_Datapath_MV2_check_n17), .ZN(
        constructing_unit_Datapath_UA_flag[2]) );
  INV_X1 constructing_unit_Datapath_UA_flag_1st_delay_U3 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_UA_flag_1st_delay_n1) );
  DFFR_X1 constructing_unit_Datapath_UA_flag_1st_delay_Q_int_reg ( .D(
        constructing_unit_Datapath_UA_flag_int_0_), .CK(clk), .RN(
        constructing_unit_Datapath_UA_flag_1st_delay_n1), .Q(
        constructing_unit_Datapath_UA_flag_int_1_) );
  INV_X1 constructing_unit_Datapath_UA_flag_delay_FFX_2_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_UA_flag_delay_FFX_2_n1) );
  DFFR_X1 constructing_unit_Datapath_UA_flag_delay_FFX_2_Q_int_reg ( .D(
        constructing_unit_Datapath_UA_flag_int_1_), .CK(clk), .RN(
        constructing_unit_Datapath_UA_flag_delay_FFX_2_n1), .Q(
        constructing_unit_Datapath_UA_flag_int_2_) );
  INV_X1 constructing_unit_Datapath_UA_flag_delay_FFX_3_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_UA_flag_delay_FFX_3_n1) );
  DFFR_X1 constructing_unit_Datapath_UA_flag_delay_FFX_3_Q_int_reg ( .D(
        constructing_unit_Datapath_UA_flag_int_2_), .CK(clk), .RN(
        constructing_unit_Datapath_UA_flag_delay_FFX_3_n1), .Q(
        constructing_unit_Datapath_UA_flag_int_3_) );
  INV_X1 constructing_unit_Datapath_UA_flag_delay_FFX_4_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_UA_flag_delay_FFX_4_n1) );
  DFFR_X1 constructing_unit_Datapath_UA_flag_delay_FFX_4_Q_int_reg ( .D(
        constructing_unit_Datapath_UA_flag_int_3_), .CK(clk), .RN(
        constructing_unit_Datapath_UA_flag_delay_FFX_4_n1), .Q(
        constructing_unit_Datapath_UA_flag_int_4_) );
  INV_X1 constructing_unit_Datapath_UA_flag_delay_FFX_5_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_UA_flag_delay_FFX_5_n1) );
  DFFR_X1 constructing_unit_Datapath_UA_flag_delay_FFX_5_Q_int_reg ( .D(
        constructing_unit_Datapath_UA_flag_int_4_), .CK(clk), .RN(
        constructing_unit_Datapath_UA_flag_delay_FFX_5_n1), .Q(
        constructing_unit_Datapath_UA_flag_int_5_) );
  INV_X1 constructing_unit_Datapath_UA_flag_delay_FFX_6_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_UA_flag_delay_FFX_6_n1) );
  DFFR_X1 constructing_unit_Datapath_UA_flag_delay_FFX_6_Q_int_reg ( .D(
        constructing_unit_Datapath_UA_flag_int_5_), .CK(clk), .RN(
        constructing_unit_Datapath_UA_flag_delay_FFX_6_n1), .Q(
        constructing_unit_Datapath_UA_flag_int_6_) );
  INV_X1 constructing_unit_Datapath_UA_flag_delay_FFX_7_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_UA_flag_delay_FFX_7_n1) );
  DFFR_X1 constructing_unit_Datapath_UA_flag_delay_FFX_7_Q_int_reg ( .D(
        constructing_unit_Datapath_UA_flag_int_6_), .CK(clk), .RN(
        constructing_unit_Datapath_UA_flag_delay_FFX_7_n1), .Q(
        constructing_unit_Datapath_UA_flag_int_7_) );
  INV_X1 constructing_unit_Datapath_UA_flag_delay_FFX_8_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_UA_flag_delay_FFX_8_n1) );
  DFFR_X1 constructing_unit_Datapath_UA_flag_delay_FFX_8_Q_int_reg ( .D(
        constructing_unit_Datapath_UA_flag_int_7_), .CK(clk), .RN(
        constructing_unit_Datapath_UA_flag_delay_FFX_8_n1), .Q(
        constructing_unit_Datapath_UA_flag_int_8_) );
  INV_X1 constructing_unit_Datapath_UA_flag_delay_FFX_9_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_UA_flag_delay_FFX_9_n1) );
  DFFR_X1 constructing_unit_Datapath_UA_flag_delay_FFX_9_Q_int_reg ( .D(
        constructing_unit_Datapath_UA_flag_int_8_), .CK(clk), .RN(
        constructing_unit_Datapath_UA_flag_delay_FFX_9_n1), .Q(
        constructing_unit_Datapath_UA_flag_int_9_) );
  INV_X1 constructing_unit_Datapath_UA_flag_delay_FFX_10_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_UA_flag_delay_FFX_10_n1) );
  DFFR_X1 constructing_unit_Datapath_UA_flag_delay_FFX_10_Q_int_reg ( .D(
        constructing_unit_Datapath_UA_flag_int_9_), .CK(clk), .RN(
        constructing_unit_Datapath_UA_flag_delay_FFX_10_n1), .Q(
        constructing_unit_Datapath_UA_flag_int_10_) );
  INV_X2 constructing_unit_Datapath_D_h_sq_sample_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_D_h_sq_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_26_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[26]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[26]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_25_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[25]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[25]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_24_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[24]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[24]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_23_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[23]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[23]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_22_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[22]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[22]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_21_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[21]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[21]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_20_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[20]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[20]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_19_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[19]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[19]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_18_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[18]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[18]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_17_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[17]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[17]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_16_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[16]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[16]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_15_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[15]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[15]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_14_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[14]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[14]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[13]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[13]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[12]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[12]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[11]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[11]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[10]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[10]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[9]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[9]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[8]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[8]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[7]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[7]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[6]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[6]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[5]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[5]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[4]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[4]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[3]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[3]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[2]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[2]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[1]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[1]) );
  DFFR_X1 constructing_unit_Datapath_D_h_sq_sample_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_D_h_sq_tmp[0]), .CK(clk), .RN(
        constructing_unit_Datapath_D_h_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_h_sq[0]) );
  INV_X1 constructing_unit_Datapath_D_v_sq_sample_U6 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_D_v_sq_sample_n4) );
  BUF_X1 constructing_unit_Datapath_D_v_sq_sample_U5 ( .A(
        constructing_unit_Datapath_D_v_sq_sample_n4), .Z(
        constructing_unit_Datapath_D_v_sq_sample_n3) );
  BUF_X1 constructing_unit_Datapath_D_v_sq_sample_U4 ( .A(
        constructing_unit_Datapath_D_v_sq_sample_n4), .Z(
        constructing_unit_Datapath_D_v_sq_sample_n2) );
  BUF_X1 constructing_unit_Datapath_D_v_sq_sample_U3 ( .A(
        constructing_unit_Datapath_D_v_sq_sample_n4), .Z(
        constructing_unit_Datapath_D_v_sq_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[0]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_v_sq[0]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[1]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_v_sq[1]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[2]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_v_sq[2]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[3]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_v_sq[3]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[4]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_v_sq[4]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[5]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_v_sq[5]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[6]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_v_sq[6]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[7]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_v_sq[7]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[8]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_v_sq[8]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[9]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_v_sq[9]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[10]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_v_sq[10]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[11]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n1), .Q(
        constructing_unit_Datapath_D_v_sq[11]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[12]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n2), .Q(
        constructing_unit_Datapath_D_v_sq[12]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[13]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n2), .Q(
        constructing_unit_Datapath_D_v_sq[13]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_14_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[14]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n2), .Q(
        constructing_unit_Datapath_D_v_sq[14]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_15_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[15]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n2), .Q(
        constructing_unit_Datapath_D_v_sq[15]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_16_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[16]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n2), .Q(
        constructing_unit_Datapath_D_v_sq[16]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_17_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[17]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n2), .Q(
        constructing_unit_Datapath_D_v_sq[17]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_18_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[18]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n2), .Q(
        constructing_unit_Datapath_D_v_sq[18]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_19_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[19]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n2), .Q(
        constructing_unit_Datapath_D_v_sq[19]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_20_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[20]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n2), .Q(
        constructing_unit_Datapath_D_v_sq[20]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_21_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[21]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n2), .Q(
        constructing_unit_Datapath_D_v_sq[21]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_22_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[22]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n2), .Q(
        constructing_unit_Datapath_D_v_sq[22]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_23_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[23]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n2), .Q(
        constructing_unit_Datapath_D_v_sq[23]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_24_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[24]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n3), .Q(
        constructing_unit_Datapath_D_v_sq[24]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_25_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[25]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n3), .Q(
        constructing_unit_Datapath_D_v_sq[25]) );
  DFFR_X1 constructing_unit_Datapath_D_v_sq_sample_Q_int_reg_26_ ( .D(
        constructing_unit_Datapath_D_v_sq_tmp[26]), .CK(clk), .RN(
        constructing_unit_Datapath_D_v_sq_sample_n3), .Q(
        constructing_unit_Datapath_D_v_sq[26]) );
  XOR2_X1 constructing_unit_Datapath_D_adder_add_19_U2 ( .A(
        constructing_unit_Datapath_D_v_sq[0]), .B(
        constructing_unit_Datapath_D_h_sq[0]), .Z(
        constructing_unit_Datapath_D_sq[0]) );
  AND2_X1 constructing_unit_Datapath_D_adder_add_19_U1 ( .A1(
        constructing_unit_Datapath_D_v_sq[0]), .A2(
        constructing_unit_Datapath_D_h_sq[0]), .ZN(
        constructing_unit_Datapath_D_adder_add_19_n1) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_1 ( .A(
        constructing_unit_Datapath_D_h_sq[1]), .B(
        constructing_unit_Datapath_D_v_sq[1]), .CI(
        constructing_unit_Datapath_D_adder_add_19_n1), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[2]), .S(
        constructing_unit_Datapath_D_sq[1]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_2 ( .A(
        constructing_unit_Datapath_D_h_sq[2]), .B(
        constructing_unit_Datapath_D_v_sq[2]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[2]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[3]), .S(
        constructing_unit_Datapath_D_sq[2]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_3 ( .A(
        constructing_unit_Datapath_D_h_sq[3]), .B(
        constructing_unit_Datapath_D_v_sq[3]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[3]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[4]), .S(
        constructing_unit_Datapath_D_sq[3]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_4 ( .A(
        constructing_unit_Datapath_D_h_sq[4]), .B(
        constructing_unit_Datapath_D_v_sq[4]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[4]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[5]), .S(
        constructing_unit_Datapath_D_sq[4]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_5 ( .A(
        constructing_unit_Datapath_D_h_sq[5]), .B(
        constructing_unit_Datapath_D_v_sq[5]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[5]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[6]), .S(
        constructing_unit_Datapath_D_sq[5]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_6 ( .A(
        constructing_unit_Datapath_D_h_sq[6]), .B(
        constructing_unit_Datapath_D_v_sq[6]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[6]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[7]), .S(
        constructing_unit_Datapath_D_sq[6]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_7 ( .A(
        constructing_unit_Datapath_D_h_sq[7]), .B(
        constructing_unit_Datapath_D_v_sq[7]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[7]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[8]), .S(
        constructing_unit_Datapath_D_sq[7]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_8 ( .A(
        constructing_unit_Datapath_D_h_sq[8]), .B(
        constructing_unit_Datapath_D_v_sq[8]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[8]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[9]), .S(
        constructing_unit_Datapath_D_sq[8]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_9 ( .A(
        constructing_unit_Datapath_D_h_sq[9]), .B(
        constructing_unit_Datapath_D_v_sq[9]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[9]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[10]), .S(
        constructing_unit_Datapath_D_sq[9]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_10 ( .A(
        constructing_unit_Datapath_D_h_sq[10]), .B(
        constructing_unit_Datapath_D_v_sq[10]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[10]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[11]), .S(
        constructing_unit_Datapath_D_sq[10]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_11 ( .A(
        constructing_unit_Datapath_D_h_sq[11]), .B(
        constructing_unit_Datapath_D_v_sq[11]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[11]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[12]), .S(
        constructing_unit_Datapath_D_sq[11]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_12 ( .A(
        constructing_unit_Datapath_D_h_sq[12]), .B(
        constructing_unit_Datapath_D_v_sq[12]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[12]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[13]), .S(
        constructing_unit_Datapath_D_sq[12]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_13 ( .A(
        constructing_unit_Datapath_D_h_sq[13]), .B(
        constructing_unit_Datapath_D_v_sq[13]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[13]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[14]), .S(
        constructing_unit_Datapath_D_sq[13]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_14 ( .A(
        constructing_unit_Datapath_D_h_sq[14]), .B(
        constructing_unit_Datapath_D_v_sq[14]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[14]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[15]), .S(
        constructing_unit_Datapath_D_sq[14]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_15 ( .A(
        constructing_unit_Datapath_D_h_sq[15]), .B(
        constructing_unit_Datapath_D_v_sq[15]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[15]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[16]), .S(
        constructing_unit_Datapath_D_sq[15]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_16 ( .A(
        constructing_unit_Datapath_D_h_sq[16]), .B(
        constructing_unit_Datapath_D_v_sq[16]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[16]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[17]), .S(
        constructing_unit_Datapath_D_sq[16]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_17 ( .A(
        constructing_unit_Datapath_D_h_sq[17]), .B(
        constructing_unit_Datapath_D_v_sq[17]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[17]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[18]), .S(
        constructing_unit_Datapath_D_sq[17]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_18 ( .A(
        constructing_unit_Datapath_D_h_sq[18]), .B(
        constructing_unit_Datapath_D_v_sq[18]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[18]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[19]), .S(
        constructing_unit_Datapath_D_sq[18]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_19 ( .A(
        constructing_unit_Datapath_D_h_sq[19]), .B(
        constructing_unit_Datapath_D_v_sq[19]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[19]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[20]), .S(
        constructing_unit_Datapath_D_sq[19]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_20 ( .A(
        constructing_unit_Datapath_D_h_sq[20]), .B(
        constructing_unit_Datapath_D_v_sq[20]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[20]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[21]), .S(
        constructing_unit_Datapath_D_sq[20]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_21 ( .A(
        constructing_unit_Datapath_D_h_sq[21]), .B(
        constructing_unit_Datapath_D_v_sq[21]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[21]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[22]), .S(
        constructing_unit_Datapath_D_sq[21]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_22 ( .A(
        constructing_unit_Datapath_D_h_sq[22]), .B(
        constructing_unit_Datapath_D_v_sq[22]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[22]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[23]), .S(
        constructing_unit_Datapath_D_sq[22]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_23 ( .A(
        constructing_unit_Datapath_D_h_sq[23]), .B(
        constructing_unit_Datapath_D_v_sq[23]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[23]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[24]), .S(
        constructing_unit_Datapath_D_sq[23]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_24 ( .A(
        constructing_unit_Datapath_D_h_sq[24]), .B(
        constructing_unit_Datapath_D_v_sq[24]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[24]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[25]), .S(
        constructing_unit_Datapath_D_sq[24]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_25 ( .A(
        constructing_unit_Datapath_D_h_sq[25]), .B(
        constructing_unit_Datapath_D_v_sq[25]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[25]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[26]), .S(
        constructing_unit_Datapath_D_sq[25]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_26 ( .A(
        constructing_unit_Datapath_D_h_sq[26]), .B(
        constructing_unit_Datapath_D_v_sq[26]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[26]), .CO(
        constructing_unit_Datapath_D_adder_add_19_carry[27]), .S(
        constructing_unit_Datapath_D_sq[26]) );
  FA_X1 constructing_unit_Datapath_D_adder_add_19_U1_27 ( .A(
        constructing_unit_Datapath_D_h_sq[26]), .B(
        constructing_unit_Datapath_D_v_sq[26]), .CI(
        constructing_unit_Datapath_D_adder_add_19_carry[27]), .S(
        constructing_unit_Datapath_D_sq[27]) );
  INV_X2 constructing_unit_Datapath_D_Cur_tmp_sample_U3 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_27_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[27]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[27]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_26_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[26]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[26]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_25_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[25]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[25]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_24_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[24]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[24]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_23_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[23]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[23]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_22_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[22]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[22]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_21_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[21]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[21]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_20_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[20]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[20]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_19_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[19]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[19]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_18_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[18]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[18]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_17_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[17]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[17]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_16_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[16]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[16]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_15_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[15]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[15]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_14_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[14]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[14]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[13]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[13]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[12]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[12]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[11]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[11]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[10]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[10]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[9]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[9]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[8]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[8]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[7]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[7]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[6]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[6]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[5]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[5]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[4]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[4]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[3]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[3]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[2]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[2]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[1]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[1]) );
  DFFR_X1 constructing_unit_Datapath_D_Cur_tmp_sample_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_D_Cur_tmp[0]), .CK(clk), .RN(
        constructing_unit_Datapath_D_Cur_tmp_sample_n1), .Q(D_Cur[0]) );
  INV_X1 constructing_unit_Datapath_D_D_register_U6 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_D_D_register_n4) );
  BUF_X1 constructing_unit_Datapath_D_D_register_U5 ( .A(
        constructing_unit_Datapath_D_D_register_n4), .Z(
        constructing_unit_Datapath_D_D_register_n3) );
  BUF_X1 constructing_unit_Datapath_D_D_register_U4 ( .A(
        constructing_unit_Datapath_D_D_register_n4), .Z(
        constructing_unit_Datapath_D_D_register_n2) );
  BUF_X1 constructing_unit_Datapath_D_D_register_U3 ( .A(
        constructing_unit_Datapath_D_D_register_n4), .Z(
        constructing_unit_Datapath_D_D_register_n1) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_0_ ( .D(D_Cur[0]), 
        .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n1), .Q(
        constructing_unit_Datapath_D_D_0_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_1_ ( .D(D_Cur[1]), 
        .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n1), .Q(
        constructing_unit_Datapath_D_D_1_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_2_ ( .D(D_Cur[2]), 
        .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n1), .Q(
        constructing_unit_Datapath_D_D_2_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_3_ ( .D(D_Cur[3]), 
        .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n1), .Q(
        constructing_unit_Datapath_D_D_3_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_4_ ( .D(D_Cur[4]), 
        .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n1), .Q(
        constructing_unit_Datapath_D_D_4_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_5_ ( .D(D_Cur[5]), 
        .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n1), .Q(
        constructing_unit_Datapath_D_D_5_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_6_ ( .D(D_Cur[6]), 
        .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n1), .Q(
        constructing_unit_Datapath_D_D_6_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_7_ ( .D(D_Cur[7]), 
        .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n1), .Q(
        constructing_unit_Datapath_D_D_7_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_8_ ( .D(D_Cur[8]), 
        .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n1), .Q(
        constructing_unit_Datapath_D_D_8_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_9_ ( .D(D_Cur[9]), 
        .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n1), .Q(
        constructing_unit_Datapath_D_D_9_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_10_ ( .D(D_Cur[10]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n1), .Q(
        constructing_unit_Datapath_D_D_10_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_11_ ( .D(D_Cur[11]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n1), .Q(
        constructing_unit_Datapath_D_D_11_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_12_ ( .D(D_Cur[12]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n2), .Q(
        constructing_unit_Datapath_D_D_12_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_13_ ( .D(D_Cur[13]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n2), .Q(
        constructing_unit_Datapath_D_D_13_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_14_ ( .D(D_Cur[14]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n2), .Q(
        constructing_unit_Datapath_D_D_14_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_15_ ( .D(D_Cur[15]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n2), .Q(
        constructing_unit_Datapath_D_D_15_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_16_ ( .D(D_Cur[16]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n2), .Q(
        constructing_unit_Datapath_D_D_16_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_17_ ( .D(D_Cur[17]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n2), .Q(
        constructing_unit_Datapath_D_D_17_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_18_ ( .D(D_Cur[18]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n2), .Q(
        constructing_unit_Datapath_D_D_18_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_19_ ( .D(D_Cur[19]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n2), .Q(
        constructing_unit_Datapath_D_D_19_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_20_ ( .D(D_Cur[20]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n2), .Q(
        constructing_unit_Datapath_D_D_20_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_21_ ( .D(D_Cur[21]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n2), .Q(
        constructing_unit_Datapath_D_D_21_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_22_ ( .D(D_Cur[22]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n2), .Q(
        constructing_unit_Datapath_D_D_22_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_23_ ( .D(D_Cur[23]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n2), .Q(
        constructing_unit_Datapath_D_D_23_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_24_ ( .D(D_Cur[24]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n3), .Q(
        constructing_unit_Datapath_D_D_24_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_25_ ( .D(D_Cur[25]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n3), .Q(
        constructing_unit_Datapath_D_D_25_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_26_ ( .D(D_Cur[26]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n3), .Q(
        constructing_unit_Datapath_D_D_26_) );
  DFFR_X1 constructing_unit_Datapath_D_D_register_Q_int_reg_27_ ( .D(D_Cur[27]), .CK(clk), .RN(constructing_unit_Datapath_D_D_register_n3), .Q(
        constructing_unit_Datapath_D_D_27_) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U65 ( .A1(
        constructing_unit_Datapath_D_D_19_), .A2(
        constructing_unit_Datapath_D_min_register_n89), .ZN(
        constructing_unit_Datapath_D_min_register_n20) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U64 ( .B1(
        constructing_unit_Datapath_D_min_register_n48), .B2(
        constructing_unit_Datapath_D_min_register_n89), .A(
        constructing_unit_Datapath_D_min_register_n20), .ZN(
        constructing_unit_Datapath_D_min_register_n76) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U63 ( .A1(
        constructing_unit_Datapath_D_D_18_), .A2(
        constructing_unit_Datapath_D_min_register_n89), .ZN(
        constructing_unit_Datapath_D_min_register_n19) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U62 ( .B1(
        constructing_unit_Datapath_D_min_register_n47), .B2(
        constructing_unit_Datapath_D_min_register_n90), .A(
        constructing_unit_Datapath_D_min_register_n19), .ZN(
        constructing_unit_Datapath_D_min_register_n75) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U61 ( .A1(
        constructing_unit_Datapath_D_D_16_), .A2(
        constructing_unit_Datapath_D_min_register_n89), .ZN(
        constructing_unit_Datapath_D_min_register_n17) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U60 ( .B1(
        constructing_unit_Datapath_D_min_register_n45), .B2(
        constructing_unit_Datapath_D_min_register_n90), .A(
        constructing_unit_Datapath_D_min_register_n17), .ZN(
        constructing_unit_Datapath_D_min_register_n73) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U59 ( .A1(
        constructing_unit_Datapath_D_D_26_), .A2(
        constructing_unit_Datapath_D_min_register_n87), .ZN(
        constructing_unit_Datapath_D_min_register_n27) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U58 ( .B1(
        constructing_unit_Datapath_D_min_register_n55), .B2(
        constructing_unit_Datapath_D_min_register_n89), .A(
        constructing_unit_Datapath_D_min_register_n27), .ZN(
        constructing_unit_Datapath_D_min_register_n83) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U57 ( .A1(
        constructing_unit_Datapath_D_D_25_), .A2(
        constructing_unit_Datapath_D_min_register_n87), .ZN(
        constructing_unit_Datapath_D_min_register_n26) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U56 ( .B1(
        constructing_unit_Datapath_D_min_register_n54), .B2(
        constructing_unit_Datapath_D_min_register_n89), .A(
        constructing_unit_Datapath_D_min_register_n26), .ZN(
        constructing_unit_Datapath_D_min_register_n82) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U55 ( .A1(
        constructing_unit_Datapath_D_D_24_), .A2(
        constructing_unit_Datapath_D_min_register_n87), .ZN(
        constructing_unit_Datapath_D_min_register_n25) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U54 ( .B1(
        constructing_unit_Datapath_D_min_register_n53), .B2(
        constructing_unit_Datapath_D_min_register_n89), .A(
        constructing_unit_Datapath_D_min_register_n25), .ZN(
        constructing_unit_Datapath_D_min_register_n81) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U53 ( .A1(
        constructing_unit_Datapath_D_D_23_), .A2(
        constructing_unit_Datapath_D_min_register_n87), .ZN(
        constructing_unit_Datapath_D_min_register_n24) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U52 ( .B1(
        constructing_unit_Datapath_D_min_register_n52), .B2(
        constructing_unit_Datapath_D_min_register_n89), .A(
        constructing_unit_Datapath_D_min_register_n24), .ZN(
        constructing_unit_Datapath_D_min_register_n80) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U51 ( .A1(
        constructing_unit_Datapath_D_D_22_), .A2(
        constructing_unit_Datapath_D_min_register_n88), .ZN(
        constructing_unit_Datapath_D_min_register_n23) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U50 ( .B1(
        constructing_unit_Datapath_D_min_register_n51), .B2(
        constructing_unit_Datapath_D_min_register_n89), .A(
        constructing_unit_Datapath_D_min_register_n23), .ZN(
        constructing_unit_Datapath_D_min_register_n79) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U49 ( .A1(
        constructing_unit_Datapath_D_D_21_), .A2(
        constructing_unit_Datapath_D_min_register_n88), .ZN(
        constructing_unit_Datapath_D_min_register_n22) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U48 ( .B1(
        constructing_unit_Datapath_D_min_register_n50), .B2(
        constructing_unit_Datapath_D_min_register_n89), .A(
        constructing_unit_Datapath_D_min_register_n22), .ZN(
        constructing_unit_Datapath_D_min_register_n78) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U47 ( .A1(
        constructing_unit_Datapath_D_D_20_), .A2(
        constructing_unit_Datapath_D_min_register_n88), .ZN(
        constructing_unit_Datapath_D_min_register_n21) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U46 ( .B1(
        constructing_unit_Datapath_D_min_register_n49), .B2(
        constructing_unit_Datapath_D_min_register_n89), .A(
        constructing_unit_Datapath_D_min_register_n21), .ZN(
        constructing_unit_Datapath_D_min_register_n77) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U45 ( .A1(
        constructing_unit_Datapath_D_D_17_), .A2(
        constructing_unit_Datapath_D_min_register_n88), .ZN(
        constructing_unit_Datapath_D_min_register_n18) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U44 ( .B1(
        constructing_unit_Datapath_D_min_register_n46), .B2(
        constructing_unit_Datapath_D_min_register_n90), .A(
        constructing_unit_Datapath_D_min_register_n18), .ZN(
        constructing_unit_Datapath_D_min_register_n74) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U43 ( .A1(
        constructing_unit_Datapath_D_D_15_), .A2(
        constructing_unit_Datapath_D_min_register_n88), .ZN(
        constructing_unit_Datapath_D_min_register_n16) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U42 ( .B1(
        constructing_unit_Datapath_D_min_register_n44), .B2(
        constructing_unit_Datapath_D_min_register_n90), .A(
        constructing_unit_Datapath_D_min_register_n16), .ZN(
        constructing_unit_Datapath_D_min_register_n72) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U41 ( .A1(
        constructing_unit_Datapath_D_D_14_), .A2(
        constructing_unit_Datapath_D_min_register_n88), .ZN(
        constructing_unit_Datapath_D_min_register_n15) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U40 ( .B1(
        constructing_unit_Datapath_D_min_register_n43), .B2(
        constructing_unit_Datapath_D_min_register_n90), .A(
        constructing_unit_Datapath_D_min_register_n15), .ZN(
        constructing_unit_Datapath_D_min_register_n71) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U39 ( .A1(
        constructing_unit_Datapath_D_D_13_), .A2(
        constructing_unit_Datapath_D_min_register_n88), .ZN(
        constructing_unit_Datapath_D_min_register_n14) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U38 ( .B1(
        constructing_unit_Datapath_D_min_register_n42), .B2(
        constructing_unit_Datapath_D_min_register_n90), .A(
        constructing_unit_Datapath_D_min_register_n14), .ZN(
        constructing_unit_Datapath_D_min_register_n70) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U37 ( .A1(
        constructing_unit_Datapath_D_D_12_), .A2(
        constructing_unit_Datapath_D_min_register_n88), .ZN(
        constructing_unit_Datapath_D_min_register_n13) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U36 ( .B1(
        constructing_unit_Datapath_D_min_register_n41), .B2(
        constructing_unit_Datapath_D_min_register_n90), .A(
        constructing_unit_Datapath_D_min_register_n13), .ZN(
        constructing_unit_Datapath_D_min_register_n69) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U35 ( .A1(
        constructing_unit_Datapath_D_D_11_), .A2(
        constructing_unit_Datapath_D_min_register_n88), .ZN(
        constructing_unit_Datapath_D_min_register_n12) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U34 ( .B1(
        constructing_unit_Datapath_D_min_register_n40), .B2(
        constructing_unit_Datapath_D_min_register_n90), .A(
        constructing_unit_Datapath_D_min_register_n12), .ZN(
        constructing_unit_Datapath_D_min_register_n68) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U33 ( .A1(
        constructing_unit_Datapath_D_D_10_), .A2(
        constructing_unit_Datapath_D_min_register_n88), .ZN(
        constructing_unit_Datapath_D_min_register_n11) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U32 ( .B1(
        constructing_unit_Datapath_D_min_register_n39), .B2(
        constructing_unit_Datapath_D_min_register_n90), .A(
        constructing_unit_Datapath_D_min_register_n11), .ZN(
        constructing_unit_Datapath_D_min_register_n67) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U31 ( .A1(
        constructing_unit_Datapath_D_D_9_), .A2(
        constructing_unit_Datapath_D_min_register_n88), .ZN(
        constructing_unit_Datapath_D_min_register_n10) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U30 ( .B1(
        constructing_unit_Datapath_D_min_register_n38), .B2(
        constructing_unit_Datapath_D_min_register_n90), .A(
        constructing_unit_Datapath_D_min_register_n10), .ZN(
        constructing_unit_Datapath_D_min_register_n66) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U29 ( .A1(
        constructing_unit_Datapath_D_D_8_), .A2(
        constructing_unit_Datapath_D_min_register_n88), .ZN(
        constructing_unit_Datapath_D_min_register_n9) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U28 ( .B1(
        constructing_unit_Datapath_D_min_register_n37), .B2(
        constructing_unit_Datapath_D_min_register_n90), .A(
        constructing_unit_Datapath_D_min_register_n9), .ZN(
        constructing_unit_Datapath_D_min_register_n65) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U27 ( .A1(
        constructing_unit_Datapath_D_min_register_n91), .A2(
        constructing_unit_Datapath_D_D_0_), .ZN(
        constructing_unit_Datapath_D_min_register_n1) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U26 ( .B1(
        constructing_unit_Datapath_D_min_register_n29), .B2(
        constructing_unit_Datapath_D_min_register_n90), .A(
        constructing_unit_Datapath_D_min_register_n1), .ZN(
        constructing_unit_Datapath_D_min_register_n57) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U25 ( .A1(
        constructing_unit_Datapath_D_D_27_), .A2(
        constructing_unit_Datapath_D_min_register_n87), .ZN(
        constructing_unit_Datapath_D_min_register_n28) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U24 ( .B1(
        constructing_unit_Datapath_D_min_register_n56), .B2(
        constructing_unit_Datapath_D_min_register_n89), .A(
        constructing_unit_Datapath_D_min_register_n28), .ZN(
        constructing_unit_Datapath_D_min_register_n85) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U23 ( .A1(
        constructing_unit_Datapath_D_D_7_), .A2(
        constructing_unit_Datapath_D_min_register_n87), .ZN(
        constructing_unit_Datapath_D_min_register_n8) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U22 ( .B1(
        constructing_unit_Datapath_D_min_register_n36), .B2(
        constructing_unit_Datapath_D_min_register_n91), .A(
        constructing_unit_Datapath_D_min_register_n8), .ZN(
        constructing_unit_Datapath_D_min_register_n64) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U21 ( .A1(
        constructing_unit_Datapath_D_D_6_), .A2(
        constructing_unit_Datapath_D_min_register_n87), .ZN(
        constructing_unit_Datapath_D_min_register_n7) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U20 ( .B1(
        constructing_unit_Datapath_D_min_register_n35), .B2(
        constructing_unit_Datapath_D_min_register_n91), .A(
        constructing_unit_Datapath_D_min_register_n7), .ZN(
        constructing_unit_Datapath_D_min_register_n63) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U19 ( .A1(
        constructing_unit_Datapath_D_D_5_), .A2(
        constructing_unit_Datapath_D_min_register_n87), .ZN(
        constructing_unit_Datapath_D_min_register_n6) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U18 ( .B1(
        constructing_unit_Datapath_D_min_register_n34), .B2(
        constructing_unit_Datapath_D_min_register_n91), .A(
        constructing_unit_Datapath_D_min_register_n6), .ZN(
        constructing_unit_Datapath_D_min_register_n62) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U17 ( .A1(
        constructing_unit_Datapath_D_D_4_), .A2(
        constructing_unit_Datapath_D_min_register_n87), .ZN(
        constructing_unit_Datapath_D_min_register_n5) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U16 ( .B1(
        constructing_unit_Datapath_D_min_register_n33), .B2(
        constructing_unit_Datapath_D_min_register_n91), .A(
        constructing_unit_Datapath_D_min_register_n5), .ZN(
        constructing_unit_Datapath_D_min_register_n61) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U15 ( .A1(
        constructing_unit_Datapath_D_D_3_), .A2(
        constructing_unit_Datapath_D_min_register_n87), .ZN(
        constructing_unit_Datapath_D_min_register_n4) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U14 ( .B1(
        constructing_unit_Datapath_D_min_register_n32), .B2(
        constructing_unit_Datapath_D_min_register_n91), .A(
        constructing_unit_Datapath_D_min_register_n4), .ZN(
        constructing_unit_Datapath_D_min_register_n60) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U13 ( .A1(
        constructing_unit_Datapath_D_D_2_), .A2(
        constructing_unit_Datapath_D_min_register_n87), .ZN(
        constructing_unit_Datapath_D_min_register_n3) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U12 ( .B1(
        constructing_unit_Datapath_D_min_register_n31), .B2(
        constructing_unit_Datapath_D_min_register_n91), .A(
        constructing_unit_Datapath_D_min_register_n3), .ZN(
        constructing_unit_Datapath_D_min_register_n59) );
  NAND2_X1 constructing_unit_Datapath_D_min_register_U11 ( .A1(
        constructing_unit_Datapath_D_D_1_), .A2(
        constructing_unit_Datapath_D_min_register_n87), .ZN(
        constructing_unit_Datapath_D_min_register_n2) );
  OAI21_X1 constructing_unit_Datapath_D_min_register_U10 ( .B1(
        constructing_unit_Datapath_D_min_register_n30), .B2(
        constructing_unit_Datapath_D_min_register_n91), .A(
        constructing_unit_Datapath_D_min_register_n2), .ZN(
        constructing_unit_Datapath_D_min_register_n58) );
  BUF_X1 constructing_unit_Datapath_D_min_register_U9 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_D_min_register_n86) );
  BUF_X1 constructing_unit_Datapath_D_min_register_U8 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_D_min_register_n84) );
  BUF_X1 constructing_unit_Datapath_D_min_register_U7 ( .A(
        constructing_unit_Datapath_D_min_register_n86), .Z(
        constructing_unit_Datapath_D_min_register_n91) );
  BUF_X1 constructing_unit_Datapath_D_min_register_U6 ( .A(
        constructing_unit_Datapath_D_min_register_n86), .Z(
        constructing_unit_Datapath_D_min_register_n90) );
  BUF_X1 constructing_unit_Datapath_D_min_register_U5 ( .A(
        constructing_unit_Datapath_D_min_register_n84), .Z(
        constructing_unit_Datapath_D_min_register_n89) );
  BUF_X1 constructing_unit_Datapath_D_min_register_U4 ( .A(
        constructing_unit_Datapath_D_min_register_n84), .Z(
        constructing_unit_Datapath_D_min_register_n87) );
  BUF_X1 constructing_unit_Datapath_D_min_register_U3 ( .A(
        constructing_unit_Datapath_D_min_register_n84), .Z(
        constructing_unit_Datapath_D_min_register_n88) );
  INV_X2 constructing_unit_Datapath_D_min_register_U2 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_D_min_register_n92) );
  DFFS_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_27_ ( .D(
        constructing_unit_Datapath_D_min_register_n85), .CK(clk), .SN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[27]), .QN(
        constructing_unit_Datapath_D_min_register_n56) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_20_ ( .D(
        constructing_unit_Datapath_D_min_register_n77), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[20]), .QN(
        constructing_unit_Datapath_D_min_register_n49) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_21_ ( .D(
        constructing_unit_Datapath_D_min_register_n78), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[21]), .QN(
        constructing_unit_Datapath_D_min_register_n50) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_22_ ( .D(
        constructing_unit_Datapath_D_min_register_n79), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[22]), .QN(
        constructing_unit_Datapath_D_min_register_n51) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_23_ ( .D(
        constructing_unit_Datapath_D_min_register_n80), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[23]), .QN(
        constructing_unit_Datapath_D_min_register_n52) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_24_ ( .D(
        constructing_unit_Datapath_D_min_register_n81), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[24]), .QN(
        constructing_unit_Datapath_D_min_register_n53) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_25_ ( .D(
        constructing_unit_Datapath_D_min_register_n82), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[25]), .QN(
        constructing_unit_Datapath_D_min_register_n54) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_26_ ( .D(
        constructing_unit_Datapath_D_min_register_n83), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[26]), .QN(
        constructing_unit_Datapath_D_min_register_n55) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_8_ ( .D(
        constructing_unit_Datapath_D_min_register_n65), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[8]), .QN(
        constructing_unit_Datapath_D_min_register_n37) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_9_ ( .D(
        constructing_unit_Datapath_D_min_register_n66), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[9]), .QN(
        constructing_unit_Datapath_D_min_register_n38) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_10_ ( .D(
        constructing_unit_Datapath_D_min_register_n67), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[10]), .QN(
        constructing_unit_Datapath_D_min_register_n39) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_11_ ( .D(
        constructing_unit_Datapath_D_min_register_n68), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[11]), .QN(
        constructing_unit_Datapath_D_min_register_n40) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_12_ ( .D(
        constructing_unit_Datapath_D_min_register_n69), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[12]), .QN(
        constructing_unit_Datapath_D_min_register_n41) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_13_ ( .D(
        constructing_unit_Datapath_D_min_register_n70), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[13]), .QN(
        constructing_unit_Datapath_D_min_register_n42) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_14_ ( .D(
        constructing_unit_Datapath_D_min_register_n71), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[14]), .QN(
        constructing_unit_Datapath_D_min_register_n43) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_15_ ( .D(
        constructing_unit_Datapath_D_min_register_n72), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[15]), .QN(
        constructing_unit_Datapath_D_min_register_n44) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_17_ ( .D(
        constructing_unit_Datapath_D_min_register_n74), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[17]), .QN(
        constructing_unit_Datapath_D_min_register_n46) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_1_ ( .D(
        constructing_unit_Datapath_D_min_register_n58), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[1]), .QN(
        constructing_unit_Datapath_D_min_register_n30) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_2_ ( .D(
        constructing_unit_Datapath_D_min_register_n59), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[2]), .QN(
        constructing_unit_Datapath_D_min_register_n31) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_3_ ( .D(
        constructing_unit_Datapath_D_min_register_n60), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[3]), .QN(
        constructing_unit_Datapath_D_min_register_n32) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_4_ ( .D(
        constructing_unit_Datapath_D_min_register_n61), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[4]), .QN(
        constructing_unit_Datapath_D_min_register_n33) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_5_ ( .D(
        constructing_unit_Datapath_D_min_register_n62), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[5]), .QN(
        constructing_unit_Datapath_D_min_register_n34) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_6_ ( .D(
        constructing_unit_Datapath_D_min_register_n63), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[6]), .QN(
        constructing_unit_Datapath_D_min_register_n35) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_7_ ( .D(
        constructing_unit_Datapath_D_min_register_n64), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[7]), .QN(
        constructing_unit_Datapath_D_min_register_n36) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_19_ ( .D(
        constructing_unit_Datapath_D_min_register_n76), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[19]), .QN(
        constructing_unit_Datapath_D_min_register_n48) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_16_ ( .D(
        constructing_unit_Datapath_D_min_register_n73), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[16]), .QN(
        constructing_unit_Datapath_D_min_register_n45) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_18_ ( .D(
        constructing_unit_Datapath_D_min_register_n75), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[18]), .QN(
        constructing_unit_Datapath_D_min_register_n47) );
  DFFR_X1 constructing_unit_Datapath_D_min_register_Q_int_reg_0_ ( .D(
        constructing_unit_Datapath_D_min_register_n57), .CK(clk), .RN(
        constructing_unit_Datapath_D_min_register_n92), .Q(
        constructing_unit_Datapath_D_min[0]), .QN(
        constructing_unit_Datapath_D_min_register_n29) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U245 ( .A1(D_Cur[9]), 
        .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n216), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n300) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U244 ( .B1(
        constructing_unit_Datapath_n68), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n233), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n300), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n304) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U243 ( .A1(D_Cur[13]), .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n213), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n294) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U242 ( .A1(D_Cur[15]), .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n212), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n296) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U241 ( .B1(
        constructing_unit_Datapath_n62), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n230), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n296), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n305) );
  OAI211_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U240 ( .C1(
        constructing_unit_Datapath_n64), .C2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n231), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n294), .B(
        constructing_unit_Datapath_final_comp_lt_gt_13_n211), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n288) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U239 ( .A1(D_Cur[11]), .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n215), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n302) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U238 ( .B1(
        constructing_unit_Datapath_n66), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n232), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n302), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n303) );
  NOR3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U237 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n304), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n288), .A3(
        constructing_unit_Datapath_final_comp_lt_gt_13_n303), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n268) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U236 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n302), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n232), .A3(
        constructing_unit_Datapath_n66), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n301) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U235 ( .B1(D_Cur[11]), .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n215), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n301), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n297) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U234 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n300), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n233), .A3(
        constructing_unit_Datapath_n68), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n299) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U233 ( .B1(D_Cur[9]), 
        .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n216), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n299), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n298) );
  OAI22_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U232 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n214), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n297), .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n297), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n298), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n289) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U231 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n296), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n230), .A3(
        constructing_unit_Datapath_n62), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n295) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U230 ( .B1(D_Cur[15]), .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n212), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n295), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n291) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U229 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n294), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n231), .A3(
        constructing_unit_Datapath_n64), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n293) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U228 ( .B1(D_Cur[13]), .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n213), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n293), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n292) );
  OAI22_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U227 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n211), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n291), .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n291), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n292), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n290) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U226 ( .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n288), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n289), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n290), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n269) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U225 ( .A1(D_Cur[3]), 
        .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n222), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n287) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U224 ( .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n236), .B2(
        constructing_unit_Datapath_n74), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n287), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n281) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U223 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n287), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n236), .A3(
        constructing_unit_Datapath_n74), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n286) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U222 ( .B1(D_Cur[3]), 
        .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n222), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n286), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n283) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U221 ( .A1(D_Cur[7]), 
        .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n219), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n278) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U220 ( .B1(
        constructing_unit_Datapath_n70), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n234), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n278), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n279) );
  AOI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U219 ( .B1(D_Cur[1]), 
        .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n224), .A(D_Cur[0]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n285) );
  AOI22_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U218 ( .A1(
        constructing_unit_Datapath_n75), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n237), .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n285), .B2(
        constructing_unit_Datapath_n76), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n284) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U217 ( .A1(D_Cur[5]), 
        .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n220), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n276) );
  OAI221_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U216 ( .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n223), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n283), .C1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n235), .C2(
        constructing_unit_Datapath_n72), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n276), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n282) );
  AOI211_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U215 ( .C1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n281), .C2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n221), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n279), .B(
        constructing_unit_Datapath_final_comp_lt_gt_13_n282), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n280) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U214 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n278), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n234), .A3(
        constructing_unit_Datapath_n70), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n277) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U213 ( .B1(D_Cur[7]), 
        .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n219), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n277), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n273) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U212 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n276), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n235), .A3(
        constructing_unit_Datapath_n72), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n275) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U211 ( .B1(D_Cur[5]), 
        .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n220), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n275), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n274) );
  OAI22_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U210 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n218), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n273), .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n273), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n274), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n272) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U209 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n217), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n272), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n270) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U208 ( .A1(D_Cur[17]), .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n210), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n256) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U207 ( .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n229), .B2(
        constructing_unit_Datapath_n60), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n256), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n271) );
  OAI221_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U206 ( .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n268), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n269), .C1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n269), .C2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n270), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n209), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n238) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U205 ( .A1(D_Cur[27]), .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n200), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n260) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U204 ( .A1(D_Cur[26]), .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n201), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n261) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U203 ( .A1(D_Cur[25]), .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n202), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n264) );
  OR2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U202 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n225), .A2(
        constructing_unit_Datapath_n24), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n267) );
  AND4_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U201 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n260), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n261), .A3(
        constructing_unit_Datapath_final_comp_lt_gt_13_n264), .A4(
        constructing_unit_Datapath_final_comp_lt_gt_13_n267), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n243) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U200 ( .A1(D_Cur[21]), .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n206), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n250) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U199 ( .A1(D_Cur[23]), .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n205), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n252) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U198 ( .B1(
        constructing_unit_Datapath_n26), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n226), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n252), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n266) );
  OAI211_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U197 ( .C1(
        constructing_unit_Datapath_n28), .C2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n227), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n250), .B(
        constructing_unit_Datapath_final_comp_lt_gt_13_n204), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n244) );
  NAND2_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U196 ( .A1(D_Cur[19]), .A2(constructing_unit_Datapath_final_comp_lt_gt_13_n208), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n258) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U195 ( .B1(
        constructing_unit_Datapath_n58), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n228), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n258), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n265) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U194 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n243), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n203), .A3(
        constructing_unit_Datapath_final_comp_lt_gt_13_n207), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n239) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U193 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n264), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n225), .A3(
        constructing_unit_Datapath_n24), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n263) );
  OAI221_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U192 ( .B1(
        D_Cur[25]), .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n202), 
        .C1(D_Cur[26]), .C2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n201), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n263), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n262) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U191 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n260), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n261), .A3(
        constructing_unit_Datapath_final_comp_lt_gt_13_n262), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n259) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U190 ( .B1(D_Cur[27]), .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n200), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n259), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n241) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U189 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n258), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n228), .A3(
        constructing_unit_Datapath_n58), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n257) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U188 ( .B1(D_Cur[19]), .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n208), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n257), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n253) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U187 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n256), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n229), .A3(
        constructing_unit_Datapath_n60), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n255) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U186 ( .B1(D_Cur[17]), .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n210), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n255), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n254) );
  OAI22_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U185 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n207), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n253), .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n253), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n254), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n245) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U184 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n252), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n226), .A3(
        constructing_unit_Datapath_n26), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n251) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U183 ( .B1(D_Cur[23]), .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n205), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n251), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n247) );
  NAND3_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U182 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n250), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n227), .A3(
        constructing_unit_Datapath_n28), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n249) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U181 ( .B1(D_Cur[21]), .B2(constructing_unit_Datapath_final_comp_lt_gt_13_n206), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n249), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n248) );
  OAI22_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U180 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n204), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n247), .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n247), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n248), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n246) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U179 ( .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n244), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n245), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n246), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n242) );
  OAI22_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U178 ( .A1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n241), .A2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n242), .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n243), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n241), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n240) );
  OAI21_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U177 ( .B1(
        constructing_unit_Datapath_final_comp_lt_gt_13_n238), .B2(
        constructing_unit_Datapath_final_comp_lt_gt_13_n239), .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n240), .ZN(
        constructing_unit_Datapath_comp_out_tmp) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U176 ( .A(
        constructing_unit_Datapath_n67), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n216) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U175 ( .A(
        constructing_unit_Datapath_n21), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n200) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U174 ( .A(
        constructing_unit_Datapath_n27), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n206) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U173 ( .A(
        constructing_unit_Datapath_n61), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n212) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U172 ( .A(
        constructing_unit_Datapath_n65), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n215) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U171 ( .A(
        constructing_unit_Datapath_n25), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n205) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U170 ( .A(
        constructing_unit_Datapath_n59), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n210) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U169 ( .A(
        constructing_unit_Datapath_n29), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n208) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U168 ( .A(
        constructing_unit_Datapath_n63), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n213) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U167 ( .A(
        constructing_unit_Datapath_n71), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n220) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U166 ( .A(
        constructing_unit_Datapath_n69), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n219) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U165 ( .A(
        constructing_unit_Datapath_n22), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n201) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U164 ( .A(
        constructing_unit_Datapath_n23), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n202) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U163 ( .A(D_Cur[24]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n225) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U162 ( .A(D_Cur[20]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n227) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U161 ( .A(D_Cur[12]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n231) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U160 ( .A(D_Cur[4]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n235) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U159 ( .A(D_Cur[22]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n226) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U158 ( .A(D_Cur[18]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n228) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U157 ( .A(D_Cur[14]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n230) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U156 ( .A(D_Cur[8]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n233) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U155 ( .A(D_Cur[10]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n232) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U154 ( .A(D_Cur[6]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n234) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U153 ( .A(D_Cur[16]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n229) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U152 ( .A(D_Cur[2]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n236) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U151 ( .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n303), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n214) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U150 ( .A(
        constructing_unit_Datapath_n73), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n222) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U149 ( .A(D_Cur[1]), 
        .ZN(constructing_unit_Datapath_final_comp_lt_gt_13_n237) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U148 ( .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n284), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n223) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U147 ( .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n280), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n217) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U146 ( .A(
        constructing_unit_Datapath_n75), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n224) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U145 ( .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n265), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n207) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U144 ( .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n266), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n204) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U143 ( .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n305), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n211) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U142 ( .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n271), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n209) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U141 ( .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n283), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n221) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U140 ( .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n279), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n218) );
  INV_X1 constructing_unit_Datapath_final_comp_lt_gt_13_U139 ( .A(
        constructing_unit_Datapath_final_comp_lt_gt_13_n244), .ZN(
        constructing_unit_Datapath_final_comp_lt_gt_13_n203) );
  INV_X1 constructing_unit_Datapath_comp_out_d_ff_U3 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_comp_out_d_ff_n1) );
  DFFR_X1 constructing_unit_Datapath_comp_out_d_ff_Q_int_reg ( .D(
        constructing_unit_Datapath_comp_out), .CK(clk), .RN(
        constructing_unit_Datapath_comp_out_d_ff_n1), .Q(
        constructing_unit_Datapath_comp_out_d) );
  INV_X1 constructing_unit_Datapath_COUNT_compEN_U9 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_COUNT_compEN_n8) );
  NOR2_X1 constructing_unit_Datapath_COUNT_compEN_U7 ( .A1(
        constructing_unit_Datapath_COUNT_compEN_n2), .A2(
        constructing_unit_Datapath_COUNT_compEN_n5), .ZN(
        constructing_unit_Datapath_COUNT_compEN_n1) );
  XOR2_X1 constructing_unit_Datapath_COUNT_compEN_U6 ( .A(
        constructing_unit_Datapath_COUNT_compEN_n1), .B(
        constructing_unit_Datapath_COUNT_compEN_n3), .Z(
        constructing_unit_Datapath_COUNT_compEN_n6) );
  NOR3_X1 constructing_unit_Datapath_COUNT_compEN_U4 ( .A1(
        constructing_unit_Datapath_COUNT_compEN_n10), .A2(
        constructing_unit_Datapath_COUNT_compEN_n4), .A3(
        constructing_unit_Datapath_COUNT_compEN_n5), .ZN(
        constructing_unit_CNT_compEN_OUT_int) );
  NAND2_X1 constructing_unit_Datapath_COUNT_compEN_U3 ( .A1(
        constructing_unit_CE_compEN_int), .A2(
        constructing_unit_Datapath_COUNT_compEN_n10), .ZN(
        constructing_unit_Datapath_COUNT_compEN_n2) );
  DFFR_X1 constructing_unit_Datapath_COUNT_compEN_count_reg_2_ ( .D(
        constructing_unit_Datapath_COUNT_compEN_n6), .CK(clk), .RN(
        constructing_unit_Datapath_COUNT_compEN_n8), .Q(
        constructing_unit_Datapath_COUNT_compEN_n3), .QN(
        constructing_unit_Datapath_COUNT_compEN_n4) );
  DFFR_X1 constructing_unit_Datapath_COUNT_compEN_count_reg_1_ ( .D(
        constructing_unit_Datapath_COUNT_compEN_n7), .CK(clk), .RN(
        constructing_unit_Datapath_COUNT_compEN_n8), .QN(
        constructing_unit_Datapath_COUNT_compEN_n5) );
  DFFR_X1 constructing_unit_Datapath_COUNT_compEN_count_reg_0_ ( .D(
        constructing_unit_Datapath_COUNT_compEN_n9), .CK(clk), .RN(
        constructing_unit_Datapath_COUNT_compEN_n8), .Q(
        constructing_unit_Datapath_COUNT_compEN_n10) );
  XOR2_X1 constructing_unit_Datapath_COUNT_compEN_U8 ( .A(
        constructing_unit_CE_compEN_int), .B(
        constructing_unit_Datapath_COUNT_compEN_n10), .Z(
        constructing_unit_Datapath_COUNT_compEN_n9) );
  XOR2_X1 constructing_unit_Datapath_COUNT_compEN_U5 ( .A(
        constructing_unit_Datapath_COUNT_compEN_n2), .B(
        constructing_unit_Datapath_COUNT_compEN_n5), .Z(
        constructing_unit_Datapath_COUNT_compEN_n7) );
  INV_X1 constructing_unit_Datapath_COUNT_STOPcompEN_U11 ( .A(
        constructing_unit_Datapath_n18), .ZN(
        constructing_unit_Datapath_COUNT_STOPcompEN_n3) );
  NAND2_X1 constructing_unit_Datapath_COUNT_STOPcompEN_U9 ( .A1(
        constructing_unit_Datapath_COUNT_STOPcompEN_n2), .A2(
        constructing_unit_Datapath_COUNT_STOPcompEN_n11), .ZN(
        constructing_unit_Datapath_COUNT_STOPcompEN_n1) );
  NOR2_X1 constructing_unit_Datapath_COUNT_STOPcompEN_U8 ( .A1(
        constructing_unit_Datapath_COUNT_STOPcompEN_n4), .A2(
        constructing_unit_Datapath_COUNT_STOPcompEN_n7), .ZN(
        constructing_unit_Datapath_COUNT_STOPcompEN_n2) );
  NOR4_X1 constructing_unit_Datapath_COUNT_STOPcompEN_U6 ( .A1(
        constructing_unit_Datapath_COUNT_STOPcompEN_n6), .A2(
        constructing_unit_Datapath_COUNT_STOPcompEN_n7), .A3(
        constructing_unit_Datapath_COUNT_STOPcompEN_n11), .A4(
        constructing_unit_Datapath_COUNT_STOPcompEN_n5), .ZN(
        constructing_unit_CNT_STOPcompEN_OUT_int) );
  NAND2_X1 constructing_unit_Datapath_COUNT_STOPcompEN_U4 ( .A1(cComp_EN), 
        .A2(constructing_unit_Datapath_COUNT_STOPcompEN_n5), .ZN(
        constructing_unit_Datapath_COUNT_STOPcompEN_n4) );
  DFFR_X1 constructing_unit_Datapath_COUNT_STOPcompEN_count_reg_3_ ( .D(
        constructing_unit_Datapath_COUNT_STOPcompEN_n8), .CK(clk), .RN(
        constructing_unit_Datapath_COUNT_STOPcompEN_n3), .QN(
        constructing_unit_Datapath_COUNT_STOPcompEN_n6) );
  DFFR_X1 constructing_unit_Datapath_COUNT_STOPcompEN_count_reg_2_ ( .D(
        constructing_unit_Datapath_COUNT_STOPcompEN_n9), .CK(clk), .RN(
        constructing_unit_Datapath_COUNT_STOPcompEN_n3), .Q(
        constructing_unit_Datapath_COUNT_STOPcompEN_n11) );
  DFFR_X1 constructing_unit_Datapath_COUNT_STOPcompEN_count_reg_1_ ( .D(
        constructing_unit_Datapath_COUNT_STOPcompEN_n10), .CK(clk), .RN(
        constructing_unit_Datapath_COUNT_STOPcompEN_n3), .QN(
        constructing_unit_Datapath_COUNT_STOPcompEN_n7) );
  DFFR_X1 constructing_unit_Datapath_COUNT_STOPcompEN_count_reg_0_ ( .D(
        constructing_unit_Datapath_COUNT_STOPcompEN_n12), .CK(clk), .RN(
        constructing_unit_Datapath_COUNT_STOPcompEN_n3), .Q(
        constructing_unit_Datapath_COUNT_STOPcompEN_n5) );
  XOR2_X1 constructing_unit_Datapath_COUNT_STOPcompEN_U10 ( .A(cComp_EN), .B(
        constructing_unit_Datapath_COUNT_STOPcompEN_n5), .Z(
        constructing_unit_Datapath_COUNT_STOPcompEN_n12) );
  XOR2_X1 constructing_unit_Datapath_COUNT_STOPcompEN_U7 ( .A(
        constructing_unit_Datapath_COUNT_STOPcompEN_n4), .B(
        constructing_unit_Datapath_COUNT_STOPcompEN_n7), .Z(
        constructing_unit_Datapath_COUNT_STOPcompEN_n10) );
  XOR2_X1 constructing_unit_Datapath_COUNT_STOPcompEN_U5 ( .A(
        constructing_unit_Datapath_COUNT_STOPcompEN_n2), .B(
        constructing_unit_Datapath_COUNT_STOPcompEN_n11), .Z(
        constructing_unit_Datapath_COUNT_STOPcompEN_n9) );
  XOR2_X1 constructing_unit_Datapath_COUNT_STOPcompEN_U3 ( .A(
        constructing_unit_Datapath_COUNT_STOPcompEN_n1), .B(
        constructing_unit_Datapath_COUNT_STOPcompEN_n6), .Z(
        constructing_unit_Datapath_COUNT_STOPcompEN_n8) );
  INV_X1 constructing_unit_Datapath_FaS_registers0_v_1_U24 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_1_n33) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_1_U23 ( .A1(cMV0_in[21]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_v_1_n11) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_1_U22 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_1_n22), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_1_n11), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_1_n34) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_1_U21 ( .A1(cMV0_in[20]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_v_1_n10) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_1_U20 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_1_n21), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_1_n10), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_1_n32) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_1_U19 ( .A1(cMV0_in[19]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_v_1_n9) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_1_U18 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_1_n20), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_1_n9), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_1_n31) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_1_U17 ( .A1(cMV0_in[18]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_v_1_n8) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_1_U16 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_1_n19), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_1_n8), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_1_n30) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_1_U15 ( .A1(cMV0_in[17]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_v_1_n7) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_1_U14 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_1_n18), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_1_n7), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_1_n29) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_1_U13 ( .A1(cMV0_in[16]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_v_1_n6) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_1_U12 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_1_n17), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_1_n6), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_1_n28) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_1_U11 ( .A1(cMV0_in[15]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_v_1_n5) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_1_U10 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_1_n16), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_1_n5), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_1_n27) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_1_U9 ( .A1(cMV0_in[14]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_v_1_n4) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_1_U8 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_1_n15), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_1_n4), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_1_n26) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_1_U7 ( .A1(cMV0_in[13]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_v_1_n3) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_1_U6 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_1_n14), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_1_n3), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_1_n25) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_1_U5 ( .A1(cMV0_in[12]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_v_1_n2) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_1_U4 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_1_n13), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_1_n2), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_1_n24) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_1_U3 ( .A1(cMV0_in[11]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_v_1_n1) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_1_U2 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_1_n12), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_1_n1), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_1_n23) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_1_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_1_n23), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_1__0_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_1_n12) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_1_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_1_n24), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_1__1_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_1_n13) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_1_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_1_n25), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_1__2_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_1_n14) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_1_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_1_n26), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_1__3_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_1_n15) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_1_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_1_n27), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_1__4_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_1_n16) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_1_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_1_n28), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_1__5_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_1_n17) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_1_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_1_n29), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_1__6_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_1_n18) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_1_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_1_n30), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_1__7_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_1_n19) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_1_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_1_n31), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_1__8_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_1_n20) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_1_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_1_n32), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_1__9_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_1_n21) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_1_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_1_n34), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_1__10_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_1_n22) );
  INV_X1 constructing_unit_Datapath_FaS_registers0_v_2_U24 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n33) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_2_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n57) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_2_U22 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_2_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_2_n57), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n35) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_2_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n67) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_2_U20 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_2_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_2_n67), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n45) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_2_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n66) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_2_U18 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_2_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_2_n66), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n44) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_2_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n58) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_2_U16 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_2_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_2_n58), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n36) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_2_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n59) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_2_U14 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_2_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_2_n59), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n37) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_2_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n60) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_2_U12 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_2_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_2_n60), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n38) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_2_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n63) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_2_U10 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_2_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_2_n63), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n41) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_2_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n64) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_2_U8 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_2_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_2_n64), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n42) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_2_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n65) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_2_U6 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_2_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_2_n65), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n43) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_2_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n61) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_2_U4 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_2_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_2_n61), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n39) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_v_2_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_v_1__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n62) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_v_2_U2 ( .B1(
        constructing_unit_Datapath_FaS_registers0_v_2_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_v_2_n62), .ZN(
        constructing_unit_Datapath_FaS_registers0_v_2_n40) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_2_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_2_n45), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_2__0_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_2_n56) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_2_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_2_n44), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_2__1_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_2_n55) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_2_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_2_n43), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_2__2_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_2_n54) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_2_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_2_n42), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_2__3_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_2_n53) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_2_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_2_n41), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_2__4_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_2_n52) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_2_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_2_n40), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_2__5_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_2_n51) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_2_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_2_n39), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_2__6_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_2_n50) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_2_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_2_n38), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_2__7_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_2_n49) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_2_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_2_n37), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_2__8_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_2_n48) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_2_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_2_n36), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_2__9_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_2_n47) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_v_2_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_v_2_n35), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_v_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_2__10_), .QN(
        constructing_unit_Datapath_FaS_registers0_v_2_n46) );
  INV_X1 constructing_unit_Datapath_FaS_registers1_v_1_U24 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_1_n33) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_1_U23 ( .A1(cMV1_in[21]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_v_1_n57) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_1_U22 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_1_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_1_n57), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_1_n35) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_1_U21 ( .A1(cMV1_in[20]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_v_1_n58) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_1_U20 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_1_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_1_n58), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_1_n36) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_1_U19 ( .A1(cMV1_in[19]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_v_1_n59) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_1_U18 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_1_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_1_n59), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_1_n37) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_1_U17 ( .A1(cMV1_in[18]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_v_1_n60) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_1_U16 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_1_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_1_n60), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_1_n38) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_1_U15 ( .A1(cMV1_in[17]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_v_1_n61) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_1_U14 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_1_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_1_n61), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_1_n39) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_1_U13 ( .A1(cMV1_in[16]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_v_1_n62) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_1_U12 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_1_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_1_n62), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_1_n40) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_1_U11 ( .A1(cMV1_in[15]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_v_1_n63) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_1_U10 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_1_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_1_n63), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_1_n41) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_1_U9 ( .A1(cMV1_in[14]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_v_1_n64) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_1_U8 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_1_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_1_n64), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_1_n42) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_1_U7 ( .A1(cMV1_in[13]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_v_1_n65) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_1_U6 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_1_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_1_n65), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_1_n43) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_1_U5 ( .A1(cMV1_in[12]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_v_1_n66) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_1_U4 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_1_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_1_n66), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_1_n44) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_1_U3 ( .A1(cMV1_in[11]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_v_1_n67) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_1_U2 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_1_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_1_n67), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_1_n45) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_1_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_1_n45), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_1__0_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_1_n56) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_1_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_1_n44), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_1__1_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_1_n55) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_1_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_1_n43), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_1__2_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_1_n54) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_1_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_1_n42), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_1__3_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_1_n53) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_1_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_1_n41), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_1__4_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_1_n52) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_1_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_1_n40), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_1__5_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_1_n51) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_1_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_1_n39), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_1__6_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_1_n50) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_1_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_1_n38), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_1__7_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_1_n49) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_1_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_1_n37), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_1__8_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_1_n48) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_1_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_1_n36), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_1__9_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_1_n47) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_1_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_1_n35), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_1__10_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_1_n46) );
  INV_X1 constructing_unit_Datapath_FaS_registers1_v_2_U24 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n33) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_2_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n66) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_2_U22 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_2_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_2_n66), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n44) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_2_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n58) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_2_U20 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_2_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_2_n58), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n36) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_2_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n59) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_2_U18 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_2_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_2_n59), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n37) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_2_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n60) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_2_U16 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_2_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_2_n60), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n38) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_2_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n63) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_2_U14 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_2_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_2_n63), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n41) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_2_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n64) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_2_U12 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_2_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_2_n64), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n42) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_2_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n65) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_2_U10 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_2_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_2_n65), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n43) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_2_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n61) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_2_U8 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_2_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_2_n61), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n39) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_2_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n62) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_2_U6 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_2_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_2_n62), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n40) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_2_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n57) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_2_U4 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_2_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_2_n57), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n35) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_v_2_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_v_1__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n67) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_v_2_U2 ( .B1(
        constructing_unit_Datapath_FaS_registers1_v_2_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_v_2_n67), .ZN(
        constructing_unit_Datapath_FaS_registers1_v_2_n45) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_2_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_2_n45), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_2__0_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_2_n56) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_2_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_2_n44), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_2__1_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_2_n55) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_2_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_2_n43), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_2__2_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_2_n54) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_2_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_2_n42), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_2__3_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_2_n53) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_2_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_2_n41), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_2__4_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_2_n52) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_2_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_2_n40), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_2__5_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_2_n51) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_2_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_2_n39), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_2__6_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_2_n50) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_2_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_2_n38), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_2__7_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_2_n49) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_2_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_2_n37), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_2__8_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_2_n48) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_2_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_2_n36), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_2__9_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_2_n47) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_v_2_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_v_2_n35), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_v_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_2__10_), .QN(
        constructing_unit_Datapath_FaS_registers1_v_2_n46) );
  INV_X1 constructing_unit_Datapath_FaS_registers2_v_1_U24 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_1_n33) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_1_U23 ( .A1(cMV2_in[21]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_v_1_n57) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_1_U22 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_1_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_1_n57), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_1_n35) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_1_U21 ( .A1(cMV2_in[20]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_v_1_n58) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_1_U20 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_1_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_1_n58), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_1_n36) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_1_U19 ( .A1(cMV2_in[19]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_v_1_n59) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_1_U18 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_1_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_1_n59), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_1_n37) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_1_U17 ( .A1(cMV2_in[18]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_v_1_n60) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_1_U16 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_1_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_1_n60), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_1_n38) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_1_U15 ( .A1(cMV2_in[17]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_v_1_n61) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_1_U14 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_1_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_1_n61), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_1_n39) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_1_U13 ( .A1(cMV2_in[16]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_v_1_n62) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_1_U12 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_1_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_1_n62), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_1_n40) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_1_U11 ( .A1(cMV2_in[15]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_v_1_n63) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_1_U10 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_1_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_1_n63), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_1_n41) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_1_U9 ( .A1(cMV2_in[14]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_v_1_n64) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_1_U8 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_1_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_1_n64), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_1_n42) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_1_U7 ( .A1(cMV2_in[13]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_v_1_n65) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_1_U6 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_1_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_1_n65), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_1_n43) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_1_U5 ( .A1(cMV2_in[12]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_v_1_n66) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_1_U4 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_1_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_1_n66), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_1_n44) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_1_U3 ( .A1(cMV2_in[11]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_v_1_n67) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_1_U2 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_1_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_1_n67), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_1_n45) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_1_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_1_n45), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_1__0_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_1_n56) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_1_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_1_n44), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_1__1_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_1_n55) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_1_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_1_n43), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_1__2_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_1_n54) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_1_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_1_n42), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_1__3_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_1_n53) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_1_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_1_n41), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_1__4_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_1_n52) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_1_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_1_n40), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_1__5_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_1_n51) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_1_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_1_n39), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_1__6_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_1_n50) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_1_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_1_n38), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_1__7_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_1_n49) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_1_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_1_n37), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_1__8_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_1_n48) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_1_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_1_n36), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_1__9_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_1_n47) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_1_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_1_n35), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_1__10_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_1_n46) );
  INV_X1 constructing_unit_Datapath_FaS_registers2_v_2_U24 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n33) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_2_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n62) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_2_U22 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_2_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_2_n62), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n40) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_2_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n57) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_2_U20 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_2_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_2_n57), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n35) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_2_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n67) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_2_U18 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_2_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_2_n67), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n45) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_2_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n66) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_2_U16 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_2_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_2_n66), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n44) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_2_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n58) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_2_U14 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_2_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_2_n58), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n36) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_2_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n59) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_2_U12 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_2_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_2_n59), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n37) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_2_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n60) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_2_U10 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_2_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_2_n60), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n38) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_2_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n63) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_2_U8 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_2_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_2_n63), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n41) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_2_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n64) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_2_U6 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_2_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_2_n64), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n42) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_2_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n65) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_2_U4 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_2_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_2_n65), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n43) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_v_2_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_v_1__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n61) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_v_2_U2 ( .B1(
        constructing_unit_Datapath_FaS_registers2_v_2_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_v_2_n61), .ZN(
        constructing_unit_Datapath_FaS_registers2_v_2_n39) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_2_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_2_n45), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_2__0_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_2_n56) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_2_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_2_n44), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_2__1_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_2_n55) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_2_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_2_n43), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_2__2_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_2_n54) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_2_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_2_n42), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_2__3_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_2_n53) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_2_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_2_n41), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_2__4_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_2_n52) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_2_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_2_n40), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_2__5_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_2_n51) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_2_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_2_n39), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_2__6_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_2_n50) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_2_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_2_n38), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_2__7_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_2_n49) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_2_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_2_n37), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_2__8_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_2_n48) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_2_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_2_n36), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_2__9_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_2_n47) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_v_2_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_v_2_n35), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_v_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_2__10_), .QN(
        constructing_unit_Datapath_FaS_registers2_v_2_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_v_3_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_3_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_v_2__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_3_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_3_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_3_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_3_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_v_2__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_3_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_3_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_3_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_3_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_v_2__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_3_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_3_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_3_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_3_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_v_2__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_3_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_3_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_3_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_3_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_v_2__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_3_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_3_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_3_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_3_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_v_2__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_3_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_3_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_3_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_3_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_2__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_3_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_3_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_3_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_3_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_v_2__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_3_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_3_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_3_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_3_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_v_2__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_3_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_3_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_3_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_3_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_v_2__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_3_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_3_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_3_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_3_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_v_2__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_3_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_3_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_3_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_3_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_3_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_3_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_3__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_3_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_3_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_3_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_3__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_3_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_3_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_3_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_3__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_3_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_3_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_3_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_3__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_3_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_3_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_3_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_3__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_3_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_3_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_3_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_3__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_3_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_3_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_3_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_3__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_3_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_3_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_3_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_3__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_3_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_3_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_3_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_3__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_3_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_3_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_3_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_3__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_3_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_3_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_3_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_3__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_3_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_v_4_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_4_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_v_3__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_4_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_4_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_4_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_4_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_v_3__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_4_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_4_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_4_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_4_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_v_3__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_4_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_4_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_4_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_4_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_v_3__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_4_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_4_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_4_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_4_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_v_3__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_4_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_4_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_4_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_4_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_v_3__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_4_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_4_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_4_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_4_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_3__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_4_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_4_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_4_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_4_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_v_3__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_4_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_4_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_4_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_4_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_v_3__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_4_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_4_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_4_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_4_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_v_3__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_4_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_4_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_4_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_4_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_v_3__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_4_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_4_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_4_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_4_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_4_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_4_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_4__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_4_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_4_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_4_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_4__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_4_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_4_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_4_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_4__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_4_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_4_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_4_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_4__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_4_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_4_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_4_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_4__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_4_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_4_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_4_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_4__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_4_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_4_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_4_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_4__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_4_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_4_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_4_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_4__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_4_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_4_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_4_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_4__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_4_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_4_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_4_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_4__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_4_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_4_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_4_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_4__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_4_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_v_5_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_5_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_v_4__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_5_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_5_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_5_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_5_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_v_4__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_5_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_5_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_5_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_5_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_v_4__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_5_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_5_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_5_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_5_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_v_4__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_5_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_5_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_5_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_5_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_v_4__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_5_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_5_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_5_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_5_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_v_4__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_5_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_5_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_5_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_5_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_4__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_5_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_5_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_5_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_5_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_v_4__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_5_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_5_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_5_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_5_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_v_4__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_5_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_5_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_5_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_5_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_v_4__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_5_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_5_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_5_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_5_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_v_4__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_5_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_5_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_5_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_5_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_5_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_5_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_5__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_5_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_5_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_5_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_5__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_5_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_5_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_5_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_5__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_5_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_5_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_5_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_5__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_5_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_5_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_5_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_5__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_5_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_5_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_5_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_5__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_5_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_5_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_5_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_5__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_5_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_5_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_5_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_5__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_5_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_5_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_5_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_5__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_5_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_5_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_5_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_5__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_5_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_5_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_5_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_5__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_5_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_v_6_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_6_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_v_5__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_6_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_6_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_6_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_6_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_v_5__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_6_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_6_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_6_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_6_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_v_5__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_6_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_6_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_6_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_6_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_v_5__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_6_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_6_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_6_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_6_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_v_5__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_6_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_6_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_6_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_6_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_v_5__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_6_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_6_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_6_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_6_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_5__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_6_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_6_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_6_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_6_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_v_5__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_6_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_6_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_6_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_6_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_v_5__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_6_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_6_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_6_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_6_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_v_5__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_6_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_6_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_6_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_6_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_v_5__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_6_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_6_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_6_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_6_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_6_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_6_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_6__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_6_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_6_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_6_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_6__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_6_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_6_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_6_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_6__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_6_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_6_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_6_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_6__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_6_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_6_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_6_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_6__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_6_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_6_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_6_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_6__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_6_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_6_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_6_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_6__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_6_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_6_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_6_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_6__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_6_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_6_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_6_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_6__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_6_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_6_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_6_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_6__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_6_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_6_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_6_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_6__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_6_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_v_7_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_7_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_v_6__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_7_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_7_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_7_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_7_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_v_6__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_7_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_7_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_7_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_7_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_v_6__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_7_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_7_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_7_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_7_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_v_6__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_7_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_7_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_7_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_7_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_v_6__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_7_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_7_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_7_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_7_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_v_6__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_7_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_7_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_7_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_7_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_6__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_7_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_7_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_7_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_7_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_v_6__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_7_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_7_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_7_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_7_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_v_6__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_7_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_7_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_7_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_7_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_v_6__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_7_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_7_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_7_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_7_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_v_6__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_7_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_7_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_7_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_7_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_7_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_7_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[0]), .QN(
        constructing_unit_Datapath_Middle_registers0_v_7_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_7_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_7_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[1]), .QN(
        constructing_unit_Datapath_Middle_registers0_v_7_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_7_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_7_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[2]), .QN(
        constructing_unit_Datapath_Middle_registers0_v_7_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_7_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_7_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[3]), .QN(
        constructing_unit_Datapath_Middle_registers0_v_7_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_7_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_7_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[4]), .QN(
        constructing_unit_Datapath_Middle_registers0_v_7_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_7_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_7_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[5]), .QN(
        constructing_unit_Datapath_Middle_registers0_v_7_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_7_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_7_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[6]), .QN(
        constructing_unit_Datapath_Middle_registers0_v_7_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_7_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_7_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[7]), .QN(
        constructing_unit_Datapath_Middle_registers0_v_7_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_7_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_7_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[8]), .QN(
        constructing_unit_Datapath_Middle_registers0_v_7_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_7_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_7_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[9]), .QN(
        constructing_unit_Datapath_Middle_registers0_v_7_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_7_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_7_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_ext[10]), .QN(
        constructing_unit_Datapath_Middle_registers0_v_7_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_v_8_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_8_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_v_ext[9]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_8_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_8_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_8_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_8_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_v_ext[8]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_8_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_8_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_8_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_8_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_v_ext[7]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_8_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_8_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_8_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_8_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_v_ext[6]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_8_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_8_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_8_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_8_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_v_ext[5]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_8_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_8_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_8_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_8_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_v_ext[4]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_8_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_8_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_8_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_8_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_ext[3]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_8_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_8_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_8_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_8_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_v_ext[2]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_8_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_8_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_8_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_8_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_v_ext[1]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_8_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_8_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_8_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_8_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_v_ext[0]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_8_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_8_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_8_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n45) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_8_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_v_ext[10]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_8_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_8_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_8_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_8_n35) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_8_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_8_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_8__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_8_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_8_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_8_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_8__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_8_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_8_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_8_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_8__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_8_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_8_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_8_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_8__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_8_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_8_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_8_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_8__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_8_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_8_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_8_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_8__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_8_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_8_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_8_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_8__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_8_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_8_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_8_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_8__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_8_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_8_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_8_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_8__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_8_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_8_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_8_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_8__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_8_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_8_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_8_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_8__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_8_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_v_9_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_9_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_v_8__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_9_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_9_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_9_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_9_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_v_8__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_9_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_9_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_9_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_9_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_v_8__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_9_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_9_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_9_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_9_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_v_8__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_9_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_9_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_9_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_9_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_v_8__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_9_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_9_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_9_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_9_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_v_8__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_9_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_9_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_9_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_9_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_8__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_9_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_9_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_9_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_9_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_v_8__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_9_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_9_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_9_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_9_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_v_8__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_9_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_9_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_9_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_9_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_v_8__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_9_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_9_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_9_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_9_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_v_8__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_9_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_9_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_9_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_9_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_9_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_9_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_9__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_9_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_9_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_9_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_9__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_9_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_9_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_9_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_9__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_9_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_9_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_9_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_9__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_9_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_9_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_9_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_9__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_9_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_9_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_9_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_9__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_9_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_9_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_9_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_9__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_9_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_9_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_9_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_9__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_9_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_9_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_9_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_9__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_9_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_9_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_9_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_9__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_9_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_9_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_9_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_9__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_9_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_v_10_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_10_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_v_9__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_10_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_10_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_10_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_10_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_v_9__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_10_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_10_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_10_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_10_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_v_9__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_10_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_10_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_10_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_10_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_v_9__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_10_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_10_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_10_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_10_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_v_9__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_10_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_10_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_10_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_10_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_v_9__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_10_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_10_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_10_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_10_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_9__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_10_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_10_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_10_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_10_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_v_9__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_10_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_10_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_10_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_10_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_v_9__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_10_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_10_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_10_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_10_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_v_9__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_10_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_10_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_10_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_10_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_v_9__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_10_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_10_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_10_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_10_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_10_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_10_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_10__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_10_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_10_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_10_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_10__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_10_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_10_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_10_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_10__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_10_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_10_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_10_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_10__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_10_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_10_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_10_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_10__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_10_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_10_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_10_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_10__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_10_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_10_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_10_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_10__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_10_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_10_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_10_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_10__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_10_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_10_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_10_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_10__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_10_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_10_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_10_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_10__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_10_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_10_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_10_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_10__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_10_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_v_11_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_11_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_v_10__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_11_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_11_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_11_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_11_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_v_10__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_11_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_11_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_11_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_11_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_v_10__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_11_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_11_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_11_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_11_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_v_10__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_11_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_11_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_11_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_11_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_v_10__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_11_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_11_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_11_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_11_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_v_10__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_11_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_11_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_11_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_11_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_10__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_11_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_11_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_11_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_11_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_v_10__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_11_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_11_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_11_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_11_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_v_10__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_11_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_11_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_11_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_11_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_v_10__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_11_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_11_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_11_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_11_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_v_10__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_11_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_11_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_11_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_11_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_11_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_11_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_11__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_11_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_11_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_11_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_11__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_11_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_11_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_11_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_11__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_11_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_11_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_11_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_11__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_11_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_11_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_11_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_11__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_11_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_11_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_11_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_11__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_11_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_11_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_11_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_11__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_11_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_11_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_11_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_11__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_11_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_11_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_11_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_11__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_11_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_11_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_11_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_11__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_11_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_11_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_11_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_11__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_11_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_v_12_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_12_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_v_11__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_12_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_12_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_12_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_12_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_v_11__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_12_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_12_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_12_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_12_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_v_11__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_12_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_12_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_12_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_12_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_v_11__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_12_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_12_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_12_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_12_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_v_11__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_12_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_12_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_12_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_12_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_v_11__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_12_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_12_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_12_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_12_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_11__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_12_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_12_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_12_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_12_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_v_11__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_12_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_12_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_12_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_12_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_v_11__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_12_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_12_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_12_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_12_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_v_11__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_12_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_12_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_12_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_12_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_v_11__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_12_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_12_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_12_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_12_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_12_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_12_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_12__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_12_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_12_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_12_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_12__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_12_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_12_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_12_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_12__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_12_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_12_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_12_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_12__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_12_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_12_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_12_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_12__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_12_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_12_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_12_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_12__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_12_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_12_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_12_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_12__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_12_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_12_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_12_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_12__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_12_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_12_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_12_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_12__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_12_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_12_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_12_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_12__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_12_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_12_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_12_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_12__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_12_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_v_13_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_13_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_v_12__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_13_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_13_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_13_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_13_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_v_12__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_13_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_13_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_13_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_13_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_v_12__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_13_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_13_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_13_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_13_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_v_12__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_13_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_13_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_13_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_13_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_v_12__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_13_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_13_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_13_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_13_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_v_12__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_13_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_13_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_13_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_13_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_12__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_13_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_13_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_13_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_13_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_v_12__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_13_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_13_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_13_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_13_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_v_12__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_13_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_13_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_13_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_13_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_v_12__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_13_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_13_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_13_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_v_13_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_v_12__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_v_13_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_v_13_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_v_13_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_v_13_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_13_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_13_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_13__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_13_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_13_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_13_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_13__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_13_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_13_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_13_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_13__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_13_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_13_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_13_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_13__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_13_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_13_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_13_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_13__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_13_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_13_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_13_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_13__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_13_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_13_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_13_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_13__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_13_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_13_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_13_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_13__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_13_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_13_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_13_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_13__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_13_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_13_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_13_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_13__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_13_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_v_13_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_v_13_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_v_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_v_13__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_v_13_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_v_3_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_3_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_v_2__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_3_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_3_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_3_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_3_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_v_2__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_3_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_3_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_3_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_3_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_v_2__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_3_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_3_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_3_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_3_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_v_2__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_3_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_3_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_3_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_3_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_v_2__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_3_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_3_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_3_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_3_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_v_2__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_3_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_3_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_3_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_3_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_2__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_3_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_3_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_3_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_3_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_v_2__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_3_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_3_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_3_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_3_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_2__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_3_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_3_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_3_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_3_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_v_2__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_3_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_3_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_3_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_3_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_v_2__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_3_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_3_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_3_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_3_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_3_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_3_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_3__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_3_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_3_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_3_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_3__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_3_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_3_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_3_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_3__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_3_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_3_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_3_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_3__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_3_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_3_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_3_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_3__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_3_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_3_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_3_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_3__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_3_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_3_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_3_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_3__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_3_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_3_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_3_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_3__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_3_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_3_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_3_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_3__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_3_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_3_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_3_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_3__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_3_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_3_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_3_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_3__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_3_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_v_4_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_4_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_v_3__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_4_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_4_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_4_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_4_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_v_3__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_4_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_4_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_4_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_4_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_v_3__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_4_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_4_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_4_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_4_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_v_3__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_4_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_4_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_4_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_4_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_v_3__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_4_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_4_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_4_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_4_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_v_3__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_4_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_4_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_4_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_4_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_3__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_4_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_4_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_4_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_4_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_v_3__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_4_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_4_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_4_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_4_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_3__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_4_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_4_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_4_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_4_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_v_3__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_4_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_4_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_4_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_4_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_v_3__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_4_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_4_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_4_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_4_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_4_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_4_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_4__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_4_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_4_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_4_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_4__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_4_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_4_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_4_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_4__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_4_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_4_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_4_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_4__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_4_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_4_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_4_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_4__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_4_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_4_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_4_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_4__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_4_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_4_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_4_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_4__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_4_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_4_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_4_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_4__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_4_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_4_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_4_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_4__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_4_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_4_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_4_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_4__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_4_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_4_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_4_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_4__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_4_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_v_5_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_5_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_v_4__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_5_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_5_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_5_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_5_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_v_4__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_5_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_5_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_5_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_5_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_v_4__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_5_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_5_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_5_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_5_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_v_4__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_5_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_5_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_5_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_5_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_v_4__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_5_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_5_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_5_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_5_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_v_4__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_5_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_5_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_5_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_5_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_4__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_5_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_5_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_5_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_5_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_v_4__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_5_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_5_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_5_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_5_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_4__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_5_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_5_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_5_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_5_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_v_4__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_5_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_5_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_5_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_5_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_v_4__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_5_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_5_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_5_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_5_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_5_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_5_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_5__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_5_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_5_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_5_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_5__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_5_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_5_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_5_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_5__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_5_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_5_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_5_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_5__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_5_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_5_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_5_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_5__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_5_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_5_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_5_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_5__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_5_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_5_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_5_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_5__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_5_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_5_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_5_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_5__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_5_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_5_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_5_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_5__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_5_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_5_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_5_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_5__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_5_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_5_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_5_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_5__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_5_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_v_6_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_6_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_v_5__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_6_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_6_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_6_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_6_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_v_5__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_6_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_6_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_6_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_6_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_v_5__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_6_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_6_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_6_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_6_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_v_5__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_6_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_6_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_6_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_6_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_v_5__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_6_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_6_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_6_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_6_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_v_5__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_6_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_6_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_6_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_6_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_5__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_6_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_6_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_6_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_6_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_v_5__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_6_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_6_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_6_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_6_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_5__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_6_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_6_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_6_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_6_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_v_5__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_6_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_6_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_6_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_6_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_v_5__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_6_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_6_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_6_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_6_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_6_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_6_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_6__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_6_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_6_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_6_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_6__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_6_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_6_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_6_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_6__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_6_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_6_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_6_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_6__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_6_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_6_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_6_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_6__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_6_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_6_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_6_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_6__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_6_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_6_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_6_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_6__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_6_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_6_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_6_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_6__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_6_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_6_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_6_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_6__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_6_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_6_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_6_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_6__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_6_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_6_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_6_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_6__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_6_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_v_7_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_7_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_v_6__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_7_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_7_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_7_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_7_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_v_6__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_7_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_7_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_7_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_7_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_v_6__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_7_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_7_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_7_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_7_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_v_6__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_7_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_7_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_7_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_7_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_v_6__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_7_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_7_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_7_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_7_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_v_6__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_7_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_7_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_7_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_7_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_6__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_7_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_7_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_7_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_7_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_v_6__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_7_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_7_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_7_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_7_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_6__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_7_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_7_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_7_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_7_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_v_6__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_7_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_7_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_7_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_7_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_v_6__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_7_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_7_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_7_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_7_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_7_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_7_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_7__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_7_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_7_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_7_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_7__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_7_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_7_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_7_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_7__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_7_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_7_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_7_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_7__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_7_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_7_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_7_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_7__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_7_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_7_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_7_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_7__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_7_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_7_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_7_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_7__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_7_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_7_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_7_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_7__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_7_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_7_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_7_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_7__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_7_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_7_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_7_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_7__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_7_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_7_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_7_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_7__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_7_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_v_8_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_8_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_v_7__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_8_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_8_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_8_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_8_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_v_7__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_8_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_8_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_8_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_8_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_v_7__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_8_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_8_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_8_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_8_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_v_7__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_8_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_8_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_8_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_8_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_v_7__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_8_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_8_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_8_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_8_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_v_7__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_8_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_8_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_8_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_8_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_7__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_8_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_8_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_8_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_8_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_v_7__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_8_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_8_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_8_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_8_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_7__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_8_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_8_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_8_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_8_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_v_7__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_8_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_8_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_8_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_8_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_v_7__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_8_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_8_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_8_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_8_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_8_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_8_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_8__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_8_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_8_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_8_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_8__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_8_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_8_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_8_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_8__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_8_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_8_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_8_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_8__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_8_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_8_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_8_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_8__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_8_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_8_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_8_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_8__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_8_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_8_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_8_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_8__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_8_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_8_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_8_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_8__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_8_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_8_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_8_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_8__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_8_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_8_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_8_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_8__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_8_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_8_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_8_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_8__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_8_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_v_9_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_9_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_v_8__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_9_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_9_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_9_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_9_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_v_8__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_9_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_9_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_9_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_9_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_v_8__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_9_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_9_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_9_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_9_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_v_8__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_9_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_9_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_9_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_9_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_v_8__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_9_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_9_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_9_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_9_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_v_8__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_9_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_9_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_9_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_9_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_8__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_9_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_9_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_9_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_9_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_v_8__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_9_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_9_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_9_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_9_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_8__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_9_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_9_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_9_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_9_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_v_8__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_9_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_9_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_9_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_9_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_v_8__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_9_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_9_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_9_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_9_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_9_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_9_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_9__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_9_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_9_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_9_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_9__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_9_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_9_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_9_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_9__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_9_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_9_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_9_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_9__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_9_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_9_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_9_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_9__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_9_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_9_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_9_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_9__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_9_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_9_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_9_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_9__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_9_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_9_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_9_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_9__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_9_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_9_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_9_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_9__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_9_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_9_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_9_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_9__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_9_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_9_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_9_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_9__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_9_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_v_10_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_10_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_v_9__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_10_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_10_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_10_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_10_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_v_9__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_10_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_10_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_10_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_10_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_v_9__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_10_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_10_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_10_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_10_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_v_9__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_10_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_10_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_10_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_10_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_v_9__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_10_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_10_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_10_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_10_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_v_9__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_10_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_10_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_10_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_10_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_9__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_10_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_10_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_10_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_10_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_v_9__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_10_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_10_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_10_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_10_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_9__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_10_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_10_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_10_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_10_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_v_9__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_10_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_10_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_10_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_10_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_v_9__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_10_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_10_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_10_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_10_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_10_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_10_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_10__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_10_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_10_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_10_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_10__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_10_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_10_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_10_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_10__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_10_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_10_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_10_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_10__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_10_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_10_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_10_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_10__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_10_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_10_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_10_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_10__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_10_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_10_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_10_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_10__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_10_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_10_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_10_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_10__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_10_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_10_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_10_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_10__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_10_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_10_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_10_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_10__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_10_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_10_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_10_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_10__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_10_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_v_11_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_11_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_v_10__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_11_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_11_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_11_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_11_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_v_10__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_11_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_11_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_11_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_11_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_v_10__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_11_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_11_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_11_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_11_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_v_10__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_11_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_11_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_11_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_11_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_v_10__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_11_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_11_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_11_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_11_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_v_10__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_11_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_11_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_11_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_11_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_10__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_11_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_11_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_11_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_11_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_v_10__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_11_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_11_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_11_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_11_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_10__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_11_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_11_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_11_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_11_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_v_10__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_11_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_11_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_11_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_11_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_v_10__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_11_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_11_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_11_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_11_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_11_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_11_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_11__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_11_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_11_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_11_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_11__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_11_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_11_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_11_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_11__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_11_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_11_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_11_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_11__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_11_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_11_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_11_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_11__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_11_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_11_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_11_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_11__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_11_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_11_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_11_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_11__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_11_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_11_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_11_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_11__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_11_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_11_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_11_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_11__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_11_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_11_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_11_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_11__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_11_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_11_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_11_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_11__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_11_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_v_12_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_12_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_v_11__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_12_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_12_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_12_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_12_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_v_11__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_12_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_12_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_12_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_12_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_v_11__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_12_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_12_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_12_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_12_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_v_11__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_12_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_12_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_12_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_12_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_v_11__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_12_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_12_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_12_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_12_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_v_11__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_12_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_12_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_12_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_12_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_11__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_12_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_12_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_12_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_12_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_v_11__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_12_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_12_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_12_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_12_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_11__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_12_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_12_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_12_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_12_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_v_11__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_12_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_12_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_12_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_12_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_v_11__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_12_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_12_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_12_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_12_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_12_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_12_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_12__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_12_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_12_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_12_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_12__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_12_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_12_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_12_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_12__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_12_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_12_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_12_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_12__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_12_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_12_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_12_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_12__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_12_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_12_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_12_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_12__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_12_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_12_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_12_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_12__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_12_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_12_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_12_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_12__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_12_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_12_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_12_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_12__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_12_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_12_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_12_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_12__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_12_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_12_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_12_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_12__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_12_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_v_13_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_13_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_v_12__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_13_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_13_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_13_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_13_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_v_12__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_13_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_13_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_13_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_13_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_v_12__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_13_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_13_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_13_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_13_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_v_12__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_13_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_13_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_13_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_13_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_v_12__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_13_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_13_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_13_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_13_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_v_12__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_13_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_13_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_13_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_13_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_12__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_13_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_13_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_13_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_13_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_v_12__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_13_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_13_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_13_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_13_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_12__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_13_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_13_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_13_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_13_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_v_12__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_13_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_13_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_13_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_v_13_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_v_12__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_v_13_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_v_13_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_v_13_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_v_13_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_13_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_13_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_13__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_13_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_13_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_13_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_13__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_13_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_13_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_13_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_13__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_13_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_13_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_13_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_13__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_13_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_13_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_13_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_13__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_13_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_13_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_13_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_13__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_13_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_13_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_13_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_13__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_13_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_13_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_13_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_13__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_13_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_13_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_13_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_13__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_13_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_13_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_13_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_13__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_13_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_v_13_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_v_13_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_v_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_v_13__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_v_13_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_v_3_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_3_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_v_2__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_3_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_3_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_3_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_3_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_v_2__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_3_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_3_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_3_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_3_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_v_2__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_3_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_3_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_3_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_3_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_v_2__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_3_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_3_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_3_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_3_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_v_2__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_3_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_3_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_3_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_3_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_v_2__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_3_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_3_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_3_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_3_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_2__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_3_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_3_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_3_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_3_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_v_2__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_3_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_3_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_3_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_3_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_v_2__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_3_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_3_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_3_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_3_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_v_2__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_3_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_3_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_3_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_3_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_v_2__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_3_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_3_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_3_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_3_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_3_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_3_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_3__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_3_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_3_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_3_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_3__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_3_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_3_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_3_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_3__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_3_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_3_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_3_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_3__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_3_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_3_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_3_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_3__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_3_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_3_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_3_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_3__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_3_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_3_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_3_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_3__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_3_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_3_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_3_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_3__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_3_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_3_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_3_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_3__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_3_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_3_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_3_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_3__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_3_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_3_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_3_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_3__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_3_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_v_4_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_4_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_v_3__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_4_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_4_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_4_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_4_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_v_3__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_4_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_4_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_4_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_4_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_v_3__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_4_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_4_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_4_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_4_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_v_3__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_4_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_4_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_4_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_4_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_v_3__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_4_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_4_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_4_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_4_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_v_3__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_4_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_4_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_4_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_4_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_3__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_4_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_4_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_4_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_4_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_v_3__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_4_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_4_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_4_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_4_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_v_3__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_4_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_4_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_4_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_4_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_v_3__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_4_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_4_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_4_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_4_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_v_3__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_4_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_4_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_4_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_4_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_4_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_4_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_4__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_4_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_4_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_4_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_4__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_4_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_4_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_4_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_4__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_4_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_4_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_4_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_4__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_4_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_4_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_4_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_4__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_4_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_4_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_4_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_4__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_4_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_4_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_4_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_4__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_4_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_4_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_4_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_4__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_4_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_4_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_4_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_4__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_4_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_4_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_4_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_4__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_4_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_4_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_4_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_4__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_4_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_v_5_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_5_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_v_4__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_5_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_5_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_5_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_5_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_v_4__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_5_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_5_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_5_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_5_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_v_4__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_5_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_5_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_5_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_5_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_v_4__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_5_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_5_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_5_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_5_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_v_4__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_5_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_5_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_5_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_5_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_v_4__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_5_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_5_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_5_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_5_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_4__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_5_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_5_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_5_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_5_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_v_4__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_5_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_5_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_5_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_5_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_v_4__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_5_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_5_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_5_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_5_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_v_4__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_5_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_5_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_5_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_5_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_v_4__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_5_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_5_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_5_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_5_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_5_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_5_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_5__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_5_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_5_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_5_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_5__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_5_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_5_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_5_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_5__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_5_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_5_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_5_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_5__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_5_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_5_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_5_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_5__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_5_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_5_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_5_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_5__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_5_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_5_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_5_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_5__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_5_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_5_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_5_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_5__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_5_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_5_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_5_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_5__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_5_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_5_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_5_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_5__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_5_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_5_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_5_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_5__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_5_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_v_6_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_6_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_v_5__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_6_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_6_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_6_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_6_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_v_5__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_6_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_6_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_6_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_6_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_v_5__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_6_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_6_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_6_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_6_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_v_5__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_6_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_6_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_6_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_6_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_v_5__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_6_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_6_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_6_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_6_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_v_5__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_6_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_6_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_6_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_6_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_5__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_6_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_6_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_6_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_6_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_v_5__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_6_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_6_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_6_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_6_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_v_5__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_6_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_6_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_6_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_6_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_v_5__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_6_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_6_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_6_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_6_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_v_5__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_6_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_6_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_6_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_6_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_6_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_6_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_6__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_6_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_6_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_6_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_6__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_6_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_6_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_6_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_6__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_6_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_6_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_6_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_6__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_6_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_6_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_6_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_6__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_6_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_6_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_6_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_6__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_6_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_6_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_6_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_6__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_6_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_6_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_6_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_6__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_6_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_6_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_6_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_6__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_6_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_6_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_6_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_6__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_6_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_6_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_6_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_6__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_6_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_v_7_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_7_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_v_6__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_7_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_7_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_7_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_7_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_v_6__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_7_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_7_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_7_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_7_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_v_6__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_7_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_7_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_7_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_7_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_v_6__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_7_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_7_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_7_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_7_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_v_6__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_7_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_7_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_7_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_7_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_v_6__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_7_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_7_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_7_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_7_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_6__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_7_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_7_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_7_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_7_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_v_6__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_7_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_7_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_7_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_7_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_v_6__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_7_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_7_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_7_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_7_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_v_6__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_7_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_7_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_7_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_7_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_v_6__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_7_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_7_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_7_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_7_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_7_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_7_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_7__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_7_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_7_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_7_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_7__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_7_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_7_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_7_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_7__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_7_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_7_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_7_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_7__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_7_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_7_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_7_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_7__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_7_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_7_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_7_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_7__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_7_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_7_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_7_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_7__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_7_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_7_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_7_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_7__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_7_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_7_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_7_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_7__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_7_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_7_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_7_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_7__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_7_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_7_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_7_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_7__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_7_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_v_8_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_8_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_v_7__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_8_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_8_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_8_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_8_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_v_7__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_8_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_8_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_8_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_8_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_v_7__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_8_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_8_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_8_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_8_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_v_7__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_8_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_8_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_8_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_8_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_v_7__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_8_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_8_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_8_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_8_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_v_7__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_8_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_8_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_8_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_8_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_7__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_8_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_8_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_8_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_8_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_v_7__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_8_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_8_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_8_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_8_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_v_7__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_8_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_8_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_8_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_8_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_v_7__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_8_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_8_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_8_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_8_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_v_7__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_8_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_8_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_8_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_8_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_8_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_8_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[0]), .QN(
        constructing_unit_Datapath_Middle_registers2_v_8_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_8_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_8_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[1]), .QN(
        constructing_unit_Datapath_Middle_registers2_v_8_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_8_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_8_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[2]), .QN(
        constructing_unit_Datapath_Middle_registers2_v_8_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_8_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_8_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[3]), .QN(
        constructing_unit_Datapath_Middle_registers2_v_8_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_8_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_8_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[4]), .QN(
        constructing_unit_Datapath_Middle_registers2_v_8_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_8_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_8_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[5]), .QN(
        constructing_unit_Datapath_Middle_registers2_v_8_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_8_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_8_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[6]), .QN(
        constructing_unit_Datapath_Middle_registers2_v_8_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_8_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_8_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[7]), .QN(
        constructing_unit_Datapath_Middle_registers2_v_8_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_8_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_8_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[8]), .QN(
        constructing_unit_Datapath_Middle_registers2_v_8_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_8_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_8_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[9]), .QN(
        constructing_unit_Datapath_Middle_registers2_v_8_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_8_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_8_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_ext[10]), .QN(
        constructing_unit_Datapath_Middle_registers2_v_8_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_v_9_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_9_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_v_ext[9]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_9_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_9_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_9_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_9_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_v_ext[8]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_9_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_9_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_9_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_9_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_v_ext[7]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_9_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_9_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_9_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_9_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_v_ext[6]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_9_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_9_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_9_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_9_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_v_ext[5]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_9_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_9_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_9_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_9_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_v_ext[4]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_9_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_9_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_9_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_9_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_ext[3]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_9_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_9_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_9_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_9_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_v_ext[2]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_9_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_9_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_9_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_9_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_v_ext[1]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_9_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_9_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_9_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_9_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_v_ext[0]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_9_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_9_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_9_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n45) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_9_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_v_ext[10]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_9_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_9_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_9_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_9_n35) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_9_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_9_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_9__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_9_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_9_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_9_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_9__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_9_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_9_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_9_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_9__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_9_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_9_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_9_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_9__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_9_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_9_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_9_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_9__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_9_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_9_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_9_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_9__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_9_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_9_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_9_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_9__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_9_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_9_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_9_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_9__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_9_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_9_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_9_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_9__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_9_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_9_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_9_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_9__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_9_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_9_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_9_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_9__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_9_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_v_10_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_10_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_v_9__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_10_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_10_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_10_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_10_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_v_9__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_10_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_10_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_10_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_10_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_v_9__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_10_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_10_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_10_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_10_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_v_9__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_10_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_10_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_10_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_10_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_v_9__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_10_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_10_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_10_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_10_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_v_9__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_10_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_10_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_10_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_10_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_9__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_10_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_10_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_10_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_10_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_v_9__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_10_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_10_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_10_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_10_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_v_9__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_10_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_10_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_10_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_10_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_v_9__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_10_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_10_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_10_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_10_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_v_9__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_10_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_10_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_10_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_10_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_10_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_10_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_10__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_10_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_10_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_10_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_10__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_10_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_10_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_10_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_10__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_10_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_10_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_10_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_10__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_10_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_10_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_10_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_10__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_10_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_10_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_10_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_10__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_10_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_10_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_10_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_10__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_10_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_10_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_10_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_10__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_10_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_10_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_10_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_10__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_10_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_10_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_10_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_10__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_10_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_10_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_10_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_10__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_10_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_v_11_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_11_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_v_10__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_11_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_11_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_11_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_11_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_v_10__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_11_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_11_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_11_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_11_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_v_10__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_11_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_11_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_11_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_11_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_v_10__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_11_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_11_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_11_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_11_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_v_10__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_11_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_11_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_11_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_11_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_v_10__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_11_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_11_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_11_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_11_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_10__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_11_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_11_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_11_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_11_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_v_10__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_11_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_11_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_11_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_11_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_v_10__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_11_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_11_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_11_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_11_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_v_10__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_11_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_11_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_11_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_11_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_v_10__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_11_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_11_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_11_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_11_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_11_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_11_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_11__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_11_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_11_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_11_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_11__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_11_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_11_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_11_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_11__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_11_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_11_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_11_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_11__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_11_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_11_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_11_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_11__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_11_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_11_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_11_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_11__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_11_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_11_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_11_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_11__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_11_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_11_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_11_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_11__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_11_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_11_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_11_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_11__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_11_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_11_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_11_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_11__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_11_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_11_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_11_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_11__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_11_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_v_12_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_12_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_v_11__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_12_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_12_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_12_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_12_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_v_11__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_12_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_12_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_12_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_12_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_v_11__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_12_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_12_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_12_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_12_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_v_11__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_12_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_12_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_12_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_12_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_v_11__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_12_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_12_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_12_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_12_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_v_11__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_12_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_12_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_12_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_12_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_11__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_12_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_12_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_12_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_12_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_v_11__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_12_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_12_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_12_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_12_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_v_11__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_12_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_12_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_12_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_12_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_v_11__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_12_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_12_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_12_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_12_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_v_11__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_12_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_12_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_12_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_12_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_12_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_12_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_12__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_12_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_12_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_12_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_12__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_12_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_12_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_12_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_12__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_12_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_12_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_12_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_12__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_12_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_12_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_12_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_12__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_12_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_12_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_12_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_12__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_12_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_12_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_12_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_12__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_12_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_12_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_12_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_12__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_12_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_12_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_12_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_12__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_12_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_12_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_12_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_12__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_12_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_12_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_12_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_12__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_12_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_v_13_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_13_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_v_12__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_13_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_13_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_13_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_13_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_v_12__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_13_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_13_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_13_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_13_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_v_12__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_13_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_13_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_13_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_13_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_v_12__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_13_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_13_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_13_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_13_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_v_12__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_13_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_13_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_13_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_13_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_v_12__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_13_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_13_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_13_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_13_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_12__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_13_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_13_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_13_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_13_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_v_12__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_13_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_13_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_13_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_13_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_v_12__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_13_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_13_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_13_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_13_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_v_12__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_13_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_13_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_13_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_v_13_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_v_12__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_v_13_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_v_13_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_v_13_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_v_13_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_13_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_13_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_13__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_13_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_13_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_13_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_13__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_13_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_13_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_13_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_13__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_13_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_13_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_13_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_13__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_13_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_13_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_13_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_13__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_13_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_13_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_13_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_13__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_13_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_13_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_13_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_13__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_13_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_13_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_13_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_13__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_13_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_13_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_13_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_13__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_13_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_13_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_13_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_13__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_13_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_v_13_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_v_13_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_v_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_v_13__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_v_13_n46) );
  INV_X1 constructing_unit_Datapath_Last_register0_v_U26 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Last_register0_v_n36) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_v_U25 ( .A1(
        constructing_unit_Datapath_MV0_int_v_13__9_), .A2(
        constructing_unit_Datapath_Last_register0_v_n33), .ZN(
        constructing_unit_Datapath_Last_register0_v_n60) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_v_U24 ( .B1(
        constructing_unit_Datapath_Last_register0_v_n49), .B2(
        constructing_unit_Datapath_Last_register0_v_n35), .A(
        constructing_unit_Datapath_Last_register0_v_n60), .ZN(
        constructing_unit_Datapath_Last_register0_v_n38) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_v_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_v_13__8_), .A2(
        constructing_unit_Datapath_Last_register0_v_n33), .ZN(
        constructing_unit_Datapath_Last_register0_v_n61) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_v_U22 ( .B1(
        constructing_unit_Datapath_Last_register0_v_n50), .B2(
        constructing_unit_Datapath_Last_register0_v_n35), .A(
        constructing_unit_Datapath_Last_register0_v_n61), .ZN(
        constructing_unit_Datapath_Last_register0_v_n39) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_v_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_v_13__7_), .A2(
        constructing_unit_Datapath_Last_register0_v_n33), .ZN(
        constructing_unit_Datapath_Last_register0_v_n62) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_v_U20 ( .B1(
        constructing_unit_Datapath_Last_register0_v_n51), .B2(
        constructing_unit_Datapath_Last_register0_v_n35), .A(
        constructing_unit_Datapath_Last_register0_v_n62), .ZN(
        constructing_unit_Datapath_Last_register0_v_n40) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_v_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_v_13__6_), .A2(
        constructing_unit_Datapath_Last_register0_v_n33), .ZN(
        constructing_unit_Datapath_Last_register0_v_n63) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_v_U18 ( .B1(
        constructing_unit_Datapath_Last_register0_v_n52), .B2(
        constructing_unit_Datapath_Last_register0_v_n35), .A(
        constructing_unit_Datapath_Last_register0_v_n63), .ZN(
        constructing_unit_Datapath_Last_register0_v_n41) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_v_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_v_13__5_), .A2(
        constructing_unit_Datapath_Last_register0_v_n33), .ZN(
        constructing_unit_Datapath_Last_register0_v_n64) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_v_U16 ( .B1(
        constructing_unit_Datapath_Last_register0_v_n53), .B2(
        constructing_unit_Datapath_Last_register0_v_n35), .A(
        constructing_unit_Datapath_Last_register0_v_n64), .ZN(
        constructing_unit_Datapath_Last_register0_v_n42) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_v_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_v_13__4_), .A2(
        constructing_unit_Datapath_Last_register0_v_n33), .ZN(
        constructing_unit_Datapath_Last_register0_v_n65) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_v_U14 ( .B1(
        constructing_unit_Datapath_Last_register0_v_n54), .B2(
        constructing_unit_Datapath_Last_register0_v_n35), .A(
        constructing_unit_Datapath_Last_register0_v_n65), .ZN(
        constructing_unit_Datapath_Last_register0_v_n43) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_v_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_v_13__3_), .A2(
        constructing_unit_Datapath_Last_register0_v_n33), .ZN(
        constructing_unit_Datapath_Last_register0_v_n66) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_v_U12 ( .B1(
        constructing_unit_Datapath_Last_register0_v_n55), .B2(
        constructing_unit_Datapath_Last_register0_v_n35), .A(
        constructing_unit_Datapath_Last_register0_v_n66), .ZN(
        constructing_unit_Datapath_Last_register0_v_n44) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_v_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_v_13__2_), .A2(
        constructing_unit_Datapath_Last_register0_v_n33), .ZN(
        constructing_unit_Datapath_Last_register0_v_n67) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_v_U10 ( .B1(
        constructing_unit_Datapath_Last_register0_v_n56), .B2(
        constructing_unit_Datapath_Last_register0_v_n35), .A(
        constructing_unit_Datapath_Last_register0_v_n67), .ZN(
        constructing_unit_Datapath_Last_register0_v_n45) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_v_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_v_13__1_), .A2(
        constructing_unit_Datapath_Last_register0_v_n33), .ZN(
        constructing_unit_Datapath_Last_register0_v_n68) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_v_U8 ( .B1(
        constructing_unit_Datapath_Last_register0_v_n57), .B2(
        constructing_unit_Datapath_Last_register0_v_n35), .A(
        constructing_unit_Datapath_Last_register0_v_n68), .ZN(
        constructing_unit_Datapath_Last_register0_v_n46) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_v_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_v_13__0_), .A2(
        constructing_unit_Datapath_Last_register0_v_n33), .ZN(
        constructing_unit_Datapath_Last_register0_v_n69) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_v_U6 ( .B1(
        constructing_unit_Datapath_Last_register0_v_n58), .B2(
        constructing_unit_Datapath_Last_register0_v_n35), .A(
        constructing_unit_Datapath_Last_register0_v_n69), .ZN(
        constructing_unit_Datapath_Last_register0_v_n47) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_v_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_v_13__10_), .A2(
        constructing_unit_Datapath_Last_register0_v_n33), .ZN(
        constructing_unit_Datapath_Last_register0_v_n59) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_v_U4 ( .B1(
        constructing_unit_Datapath_Last_register0_v_n48), .B2(
        constructing_unit_Datapath_Last_register0_v_n33), .A(
        constructing_unit_Datapath_Last_register0_v_n59), .ZN(
        constructing_unit_Datapath_Last_register0_v_n37) );
  BUF_X1 constructing_unit_Datapath_Last_register0_v_U3 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_Last_register0_v_n35) );
  BUF_X1 constructing_unit_Datapath_Last_register0_v_U2 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_Last_register0_v_n33) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_v_MV_out_int_reg_0_ ( .D(
        constructing_unit_Datapath_Last_register0_v_n47), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_v_n36), .Q(MVP0[11]), .QN(
        constructing_unit_Datapath_Last_register0_v_n58) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_v_MV_out_int_reg_1_ ( .D(
        constructing_unit_Datapath_Last_register0_v_n46), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_v_n36), .Q(MVP0[12]), .QN(
        constructing_unit_Datapath_Last_register0_v_n57) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_v_MV_out_int_reg_2_ ( .D(
        constructing_unit_Datapath_Last_register0_v_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_v_n36), .Q(MVP0[13]), .QN(
        constructing_unit_Datapath_Last_register0_v_n56) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_v_MV_out_int_reg_3_ ( .D(
        constructing_unit_Datapath_Last_register0_v_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_v_n36), .Q(MVP0[14]), .QN(
        constructing_unit_Datapath_Last_register0_v_n55) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_v_MV_out_int_reg_4_ ( .D(
        constructing_unit_Datapath_Last_register0_v_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_v_n36), .Q(MVP0[15]), .QN(
        constructing_unit_Datapath_Last_register0_v_n54) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_v_MV_out_int_reg_5_ ( .D(
        constructing_unit_Datapath_Last_register0_v_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_v_n36), .Q(MVP0[16]), .QN(
        constructing_unit_Datapath_Last_register0_v_n53) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_v_MV_out_int_reg_6_ ( .D(
        constructing_unit_Datapath_Last_register0_v_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_v_n36), .Q(MVP0[17]), .QN(
        constructing_unit_Datapath_Last_register0_v_n52) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_v_MV_out_int_reg_7_ ( .D(
        constructing_unit_Datapath_Last_register0_v_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_v_n36), .Q(MVP0[18]), .QN(
        constructing_unit_Datapath_Last_register0_v_n51) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_v_MV_out_int_reg_8_ ( .D(
        constructing_unit_Datapath_Last_register0_v_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_v_n36), .Q(MVP0[19]), .QN(
        constructing_unit_Datapath_Last_register0_v_n50) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_v_MV_out_int_reg_9_ ( .D(
        constructing_unit_Datapath_Last_register0_v_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_v_n36), .Q(MVP0[20]), .QN(
        constructing_unit_Datapath_Last_register0_v_n49) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_v_MV_out_int_reg_10_ ( .D(
        constructing_unit_Datapath_Last_register0_v_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_v_n36), .Q(MVP0[21]), .QN(
        constructing_unit_Datapath_Last_register0_v_n48) );
  INV_X1 constructing_unit_Datapath_Last_register1_v_U26 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Last_register1_v_n36) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_v_U25 ( .A1(
        constructing_unit_Datapath_MV1_int_v_13__9_), .A2(
        constructing_unit_Datapath_Last_register1_v_n33), .ZN(
        constructing_unit_Datapath_Last_register1_v_n60) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_v_U24 ( .B1(
        constructing_unit_Datapath_Last_register1_v_n49), .B2(
        constructing_unit_Datapath_Last_register1_v_n35), .A(
        constructing_unit_Datapath_Last_register1_v_n60), .ZN(
        constructing_unit_Datapath_Last_register1_v_n38) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_v_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_v_13__8_), .A2(
        constructing_unit_Datapath_Last_register1_v_n33), .ZN(
        constructing_unit_Datapath_Last_register1_v_n61) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_v_U22 ( .B1(
        constructing_unit_Datapath_Last_register1_v_n50), .B2(
        constructing_unit_Datapath_Last_register1_v_n35), .A(
        constructing_unit_Datapath_Last_register1_v_n61), .ZN(
        constructing_unit_Datapath_Last_register1_v_n39) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_v_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_v_13__7_), .A2(
        constructing_unit_Datapath_Last_register1_v_n33), .ZN(
        constructing_unit_Datapath_Last_register1_v_n62) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_v_U20 ( .B1(
        constructing_unit_Datapath_Last_register1_v_n51), .B2(
        constructing_unit_Datapath_Last_register1_v_n35), .A(
        constructing_unit_Datapath_Last_register1_v_n62), .ZN(
        constructing_unit_Datapath_Last_register1_v_n40) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_v_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_v_13__6_), .A2(
        constructing_unit_Datapath_Last_register1_v_n33), .ZN(
        constructing_unit_Datapath_Last_register1_v_n63) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_v_U18 ( .B1(
        constructing_unit_Datapath_Last_register1_v_n52), .B2(
        constructing_unit_Datapath_Last_register1_v_n35), .A(
        constructing_unit_Datapath_Last_register1_v_n63), .ZN(
        constructing_unit_Datapath_Last_register1_v_n41) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_v_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_v_13__5_), .A2(
        constructing_unit_Datapath_Last_register1_v_n33), .ZN(
        constructing_unit_Datapath_Last_register1_v_n64) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_v_U16 ( .B1(
        constructing_unit_Datapath_Last_register1_v_n53), .B2(
        constructing_unit_Datapath_Last_register1_v_n35), .A(
        constructing_unit_Datapath_Last_register1_v_n64), .ZN(
        constructing_unit_Datapath_Last_register1_v_n42) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_v_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_v_13__4_), .A2(
        constructing_unit_Datapath_Last_register1_v_n33), .ZN(
        constructing_unit_Datapath_Last_register1_v_n65) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_v_U14 ( .B1(
        constructing_unit_Datapath_Last_register1_v_n54), .B2(
        constructing_unit_Datapath_Last_register1_v_n35), .A(
        constructing_unit_Datapath_Last_register1_v_n65), .ZN(
        constructing_unit_Datapath_Last_register1_v_n43) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_v_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_v_13__3_), .A2(
        constructing_unit_Datapath_Last_register1_v_n33), .ZN(
        constructing_unit_Datapath_Last_register1_v_n66) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_v_U12 ( .B1(
        constructing_unit_Datapath_Last_register1_v_n55), .B2(
        constructing_unit_Datapath_Last_register1_v_n35), .A(
        constructing_unit_Datapath_Last_register1_v_n66), .ZN(
        constructing_unit_Datapath_Last_register1_v_n44) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_v_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_v_13__2_), .A2(
        constructing_unit_Datapath_Last_register1_v_n33), .ZN(
        constructing_unit_Datapath_Last_register1_v_n67) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_v_U10 ( .B1(
        constructing_unit_Datapath_Last_register1_v_n56), .B2(
        constructing_unit_Datapath_Last_register1_v_n35), .A(
        constructing_unit_Datapath_Last_register1_v_n67), .ZN(
        constructing_unit_Datapath_Last_register1_v_n45) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_v_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_v_13__1_), .A2(
        constructing_unit_Datapath_Last_register1_v_n33), .ZN(
        constructing_unit_Datapath_Last_register1_v_n68) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_v_U8 ( .B1(
        constructing_unit_Datapath_Last_register1_v_n57), .B2(
        constructing_unit_Datapath_Last_register1_v_n35), .A(
        constructing_unit_Datapath_Last_register1_v_n68), .ZN(
        constructing_unit_Datapath_Last_register1_v_n46) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_v_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_v_13__0_), .A2(
        constructing_unit_Datapath_Last_register1_v_n33), .ZN(
        constructing_unit_Datapath_Last_register1_v_n69) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_v_U6 ( .B1(
        constructing_unit_Datapath_Last_register1_v_n58), .B2(
        constructing_unit_Datapath_Last_register1_v_n35), .A(
        constructing_unit_Datapath_Last_register1_v_n69), .ZN(
        constructing_unit_Datapath_Last_register1_v_n47) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_v_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_v_13__10_), .A2(
        constructing_unit_Datapath_Last_register1_v_n33), .ZN(
        constructing_unit_Datapath_Last_register1_v_n59) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_v_U4 ( .B1(
        constructing_unit_Datapath_Last_register1_v_n48), .B2(
        constructing_unit_Datapath_Last_register1_v_n33), .A(
        constructing_unit_Datapath_Last_register1_v_n59), .ZN(
        constructing_unit_Datapath_Last_register1_v_n37) );
  BUF_X1 constructing_unit_Datapath_Last_register1_v_U3 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_Last_register1_v_n35) );
  BUF_X1 constructing_unit_Datapath_Last_register1_v_U2 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_Last_register1_v_n33) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_v_MV_out_int_reg_0_ ( .D(
        constructing_unit_Datapath_Last_register1_v_n47), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_v_n36), .Q(MVP1[11]), .QN(
        constructing_unit_Datapath_Last_register1_v_n58) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_v_MV_out_int_reg_1_ ( .D(
        constructing_unit_Datapath_Last_register1_v_n46), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_v_n36), .Q(MVP1[12]), .QN(
        constructing_unit_Datapath_Last_register1_v_n57) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_v_MV_out_int_reg_2_ ( .D(
        constructing_unit_Datapath_Last_register1_v_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_v_n36), .Q(MVP1[13]), .QN(
        constructing_unit_Datapath_Last_register1_v_n56) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_v_MV_out_int_reg_3_ ( .D(
        constructing_unit_Datapath_Last_register1_v_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_v_n36), .Q(MVP1[14]), .QN(
        constructing_unit_Datapath_Last_register1_v_n55) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_v_MV_out_int_reg_4_ ( .D(
        constructing_unit_Datapath_Last_register1_v_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_v_n36), .Q(MVP1[15]), .QN(
        constructing_unit_Datapath_Last_register1_v_n54) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_v_MV_out_int_reg_5_ ( .D(
        constructing_unit_Datapath_Last_register1_v_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_v_n36), .Q(MVP1[16]), .QN(
        constructing_unit_Datapath_Last_register1_v_n53) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_v_MV_out_int_reg_6_ ( .D(
        constructing_unit_Datapath_Last_register1_v_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_v_n36), .Q(MVP1[17]), .QN(
        constructing_unit_Datapath_Last_register1_v_n52) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_v_MV_out_int_reg_7_ ( .D(
        constructing_unit_Datapath_Last_register1_v_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_v_n36), .Q(MVP1[18]), .QN(
        constructing_unit_Datapath_Last_register1_v_n51) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_v_MV_out_int_reg_8_ ( .D(
        constructing_unit_Datapath_Last_register1_v_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_v_n36), .Q(MVP1[19]), .QN(
        constructing_unit_Datapath_Last_register1_v_n50) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_v_MV_out_int_reg_9_ ( .D(
        constructing_unit_Datapath_Last_register1_v_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_v_n36), .Q(MVP1[20]), .QN(
        constructing_unit_Datapath_Last_register1_v_n49) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_v_MV_out_int_reg_10_ ( .D(
        constructing_unit_Datapath_Last_register1_v_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_v_n36), .Q(MVP1[21]), .QN(
        constructing_unit_Datapath_Last_register1_v_n48) );
  INV_X1 constructing_unit_Datapath_Last_register2_v_U26 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Last_register2_v_n36) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_v_U25 ( .A1(
        constructing_unit_Datapath_MV2_int_v_13__9_), .A2(
        constructing_unit_Datapath_Last_register2_v_n33), .ZN(
        constructing_unit_Datapath_Last_register2_v_n60) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_v_U24 ( .B1(
        constructing_unit_Datapath_Last_register2_v_n49), .B2(
        constructing_unit_Datapath_Last_register2_v_n35), .A(
        constructing_unit_Datapath_Last_register2_v_n60), .ZN(
        constructing_unit_Datapath_Last_register2_v_n38) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_v_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_v_13__8_), .A2(
        constructing_unit_Datapath_Last_register2_v_n33), .ZN(
        constructing_unit_Datapath_Last_register2_v_n61) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_v_U22 ( .B1(
        constructing_unit_Datapath_Last_register2_v_n50), .B2(
        constructing_unit_Datapath_Last_register2_v_n35), .A(
        constructing_unit_Datapath_Last_register2_v_n61), .ZN(
        constructing_unit_Datapath_Last_register2_v_n39) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_v_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_v_13__7_), .A2(
        constructing_unit_Datapath_Last_register2_v_n33), .ZN(
        constructing_unit_Datapath_Last_register2_v_n62) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_v_U20 ( .B1(
        constructing_unit_Datapath_Last_register2_v_n51), .B2(
        constructing_unit_Datapath_Last_register2_v_n35), .A(
        constructing_unit_Datapath_Last_register2_v_n62), .ZN(
        constructing_unit_Datapath_Last_register2_v_n40) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_v_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_v_13__6_), .A2(
        constructing_unit_Datapath_Last_register2_v_n33), .ZN(
        constructing_unit_Datapath_Last_register2_v_n63) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_v_U18 ( .B1(
        constructing_unit_Datapath_Last_register2_v_n52), .B2(
        constructing_unit_Datapath_Last_register2_v_n35), .A(
        constructing_unit_Datapath_Last_register2_v_n63), .ZN(
        constructing_unit_Datapath_Last_register2_v_n41) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_v_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_v_13__5_), .A2(
        constructing_unit_Datapath_Last_register2_v_n33), .ZN(
        constructing_unit_Datapath_Last_register2_v_n64) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_v_U16 ( .B1(
        constructing_unit_Datapath_Last_register2_v_n53), .B2(
        constructing_unit_Datapath_Last_register2_v_n35), .A(
        constructing_unit_Datapath_Last_register2_v_n64), .ZN(
        constructing_unit_Datapath_Last_register2_v_n42) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_v_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_v_13__4_), .A2(
        constructing_unit_Datapath_Last_register2_v_n33), .ZN(
        constructing_unit_Datapath_Last_register2_v_n65) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_v_U14 ( .B1(
        constructing_unit_Datapath_Last_register2_v_n54), .B2(
        constructing_unit_Datapath_Last_register2_v_n35), .A(
        constructing_unit_Datapath_Last_register2_v_n65), .ZN(
        constructing_unit_Datapath_Last_register2_v_n43) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_v_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_v_13__3_), .A2(
        constructing_unit_Datapath_Last_register2_v_n33), .ZN(
        constructing_unit_Datapath_Last_register2_v_n66) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_v_U12 ( .B1(
        constructing_unit_Datapath_Last_register2_v_n55), .B2(
        constructing_unit_Datapath_Last_register2_v_n35), .A(
        constructing_unit_Datapath_Last_register2_v_n66), .ZN(
        constructing_unit_Datapath_Last_register2_v_n44) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_v_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_v_13__2_), .A2(
        constructing_unit_Datapath_Last_register2_v_n33), .ZN(
        constructing_unit_Datapath_Last_register2_v_n67) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_v_U10 ( .B1(
        constructing_unit_Datapath_Last_register2_v_n56), .B2(
        constructing_unit_Datapath_Last_register2_v_n35), .A(
        constructing_unit_Datapath_Last_register2_v_n67), .ZN(
        constructing_unit_Datapath_Last_register2_v_n45) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_v_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_v_13__1_), .A2(
        constructing_unit_Datapath_Last_register2_v_n33), .ZN(
        constructing_unit_Datapath_Last_register2_v_n68) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_v_U8 ( .B1(
        constructing_unit_Datapath_Last_register2_v_n57), .B2(
        constructing_unit_Datapath_Last_register2_v_n35), .A(
        constructing_unit_Datapath_Last_register2_v_n68), .ZN(
        constructing_unit_Datapath_Last_register2_v_n46) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_v_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_v_13__0_), .A2(
        constructing_unit_Datapath_Last_register2_v_n33), .ZN(
        constructing_unit_Datapath_Last_register2_v_n69) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_v_U6 ( .B1(
        constructing_unit_Datapath_Last_register2_v_n58), .B2(
        constructing_unit_Datapath_Last_register2_v_n35), .A(
        constructing_unit_Datapath_Last_register2_v_n69), .ZN(
        constructing_unit_Datapath_Last_register2_v_n47) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_v_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_v_13__10_), .A2(
        constructing_unit_Datapath_Last_register2_v_n33), .ZN(
        constructing_unit_Datapath_Last_register2_v_n59) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_v_U4 ( .B1(
        constructing_unit_Datapath_Last_register2_v_n48), .B2(
        constructing_unit_Datapath_Last_register2_v_n33), .A(
        constructing_unit_Datapath_Last_register2_v_n59), .ZN(
        constructing_unit_Datapath_Last_register2_v_n37) );
  BUF_X1 constructing_unit_Datapath_Last_register2_v_U3 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_Last_register2_v_n35) );
  BUF_X1 constructing_unit_Datapath_Last_register2_v_U2 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_Last_register2_v_n33) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_v_MV_out_int_reg_0_ ( .D(
        constructing_unit_Datapath_Last_register2_v_n47), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_v_n36), .Q(MVP2[11]), .QN(
        constructing_unit_Datapath_Last_register2_v_n58) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_v_MV_out_int_reg_1_ ( .D(
        constructing_unit_Datapath_Last_register2_v_n46), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_v_n36), .Q(MVP2[12]), .QN(
        constructing_unit_Datapath_Last_register2_v_n57) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_v_MV_out_int_reg_2_ ( .D(
        constructing_unit_Datapath_Last_register2_v_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_v_n36), .Q(MVP2[13]), .QN(
        constructing_unit_Datapath_Last_register2_v_n56) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_v_MV_out_int_reg_3_ ( .D(
        constructing_unit_Datapath_Last_register2_v_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_v_n36), .Q(MVP2[14]), .QN(
        constructing_unit_Datapath_Last_register2_v_n55) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_v_MV_out_int_reg_4_ ( .D(
        constructing_unit_Datapath_Last_register2_v_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_v_n36), .Q(MVP2[15]), .QN(
        constructing_unit_Datapath_Last_register2_v_n54) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_v_MV_out_int_reg_5_ ( .D(
        constructing_unit_Datapath_Last_register2_v_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_v_n36), .Q(MVP2[16]), .QN(
        constructing_unit_Datapath_Last_register2_v_n53) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_v_MV_out_int_reg_6_ ( .D(
        constructing_unit_Datapath_Last_register2_v_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_v_n36), .Q(MVP2[17]), .QN(
        constructing_unit_Datapath_Last_register2_v_n52) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_v_MV_out_int_reg_7_ ( .D(
        constructing_unit_Datapath_Last_register2_v_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_v_n36), .Q(MVP2[18]), .QN(
        constructing_unit_Datapath_Last_register2_v_n51) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_v_MV_out_int_reg_8_ ( .D(
        constructing_unit_Datapath_Last_register2_v_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_v_n36), .Q(MVP2[19]), .QN(
        constructing_unit_Datapath_Last_register2_v_n50) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_v_MV_out_int_reg_9_ ( .D(
        constructing_unit_Datapath_Last_register2_v_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_v_n36), .Q(MVP2[20]), .QN(
        constructing_unit_Datapath_Last_register2_v_n49) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_v_MV_out_int_reg_10_ ( .D(
        constructing_unit_Datapath_Last_register2_v_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_v_n36), .Q(MVP2[21]), .QN(
        constructing_unit_Datapath_Last_register2_v_n48) );
  INV_X1 constructing_unit_Datapath_FaS_registers0_h_1_U24 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_1_n33) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_1_U23 ( .A1(cMV0_in[10]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_h_1_n57) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_1_U22 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_1_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_1_n57), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_1_n35) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_1_U21 ( .A1(cMV0_in[9]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_h_1_n58) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_1_U20 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_1_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_1_n58), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_1_n36) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_1_U19 ( .A1(cMV0_in[8]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_h_1_n59) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_1_U18 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_1_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_1_n59), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_1_n37) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_1_U17 ( .A1(cMV0_in[7]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_h_1_n60) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_1_U16 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_1_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_1_n60), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_1_n38) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_1_U15 ( .A1(cMV0_in[6]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_h_1_n61) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_1_U14 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_1_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_1_n61), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_1_n39) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_1_U13 ( .A1(cMV0_in[5]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_h_1_n62) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_1_U12 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_1_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_1_n62), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_1_n40) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_1_U11 ( .A1(cMV0_in[4]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_h_1_n63) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_1_U10 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_1_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_1_n63), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_1_n41) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_1_U9 ( .A1(cMV0_in[3]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_h_1_n64) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_1_U8 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_1_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_1_n64), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_1_n42) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_1_U7 ( .A1(cMV0_in[2]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_h_1_n65) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_1_U6 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_1_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_1_n65), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_1_n43) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_1_U5 ( .A1(cMV0_in[1]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_h_1_n66) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_1_U4 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_1_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_1_n66), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_1_n44) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_1_U3 ( .A1(cMV0_in[0]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers0_h_1_n67) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_1_U2 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_1_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_1_n67), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_1_n45) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_1_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_1_n45), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_1__0_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_1_n56) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_1_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_1_n44), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_1__1_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_1_n55) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_1_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_1_n43), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_1__2_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_1_n54) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_1_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_1_n42), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_1__3_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_1_n53) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_1_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_1_n41), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_1__4_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_1_n52) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_1_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_1_n40), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_1__5_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_1_n51) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_1_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_1_n39), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_1__6_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_1_n50) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_1_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_1_n38), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_1__7_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_1_n49) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_1_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_1_n37), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_1__8_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_1_n48) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_1_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_1_n36), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_1__9_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_1_n47) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_1_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_1_n35), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_1_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_1__10_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_1_n46) );
  INV_X1 constructing_unit_Datapath_FaS_registers0_h_2_U24 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n33) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_2_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n57) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_2_U22 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_2_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_2_n57), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n35) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_2_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n67) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_2_U20 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_2_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_2_n67), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n45) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_2_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n66) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_2_U18 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_2_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_2_n66), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n44) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_2_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n58) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_2_U16 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_2_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_2_n58), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n36) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_2_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n59) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_2_U14 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_2_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_2_n59), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n37) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_2_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n60) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_2_U12 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_2_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_2_n60), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n38) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_2_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n63) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_2_U10 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_2_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_2_n63), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n41) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_2_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n64) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_2_U8 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_2_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_2_n64), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n42) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_2_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n65) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_2_U6 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_2_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_2_n65), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n43) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_2_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n61) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_2_U4 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_2_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_2_n61), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n39) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers0_h_2_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_h_1__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n62) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers0_h_2_U2 ( .B1(
        constructing_unit_Datapath_FaS_registers0_h_2_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers0_h_2_n62), .ZN(
        constructing_unit_Datapath_FaS_registers0_h_2_n40) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_2_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_2_n45), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_2__0_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_2_n56) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_2_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_2_n44), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_2__1_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_2_n55) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_2_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_2_n43), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_2__2_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_2_n54) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_2_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_2_n42), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_2__3_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_2_n53) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_2_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_2_n41), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_2__4_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_2_n52) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_2_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_2_n40), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_2__5_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_2_n51) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_2_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_2_n39), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_2__6_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_2_n50) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_2_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_2_n38), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_2__7_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_2_n49) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_2_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_2_n37), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_2__8_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_2_n48) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_2_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_2_n36), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_2__9_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_2_n47) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers0_h_2_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_FaS_registers0_h_2_n35), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers0_h_2_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_2__10_), .QN(
        constructing_unit_Datapath_FaS_registers0_h_2_n46) );
  INV_X1 constructing_unit_Datapath_FaS_registers1_h_1_U24 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_1_n33) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_1_U23 ( .A1(cMV1_in[10]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_h_1_n57) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_1_U22 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_1_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_1_n57), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_1_n35) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_1_U21 ( .A1(cMV1_in[9]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_h_1_n58) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_1_U20 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_1_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_1_n58), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_1_n36) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_1_U19 ( .A1(cMV1_in[8]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_h_1_n59) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_1_U18 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_1_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_1_n59), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_1_n37) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_1_U17 ( .A1(cMV1_in[7]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_h_1_n60) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_1_U16 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_1_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_1_n60), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_1_n38) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_1_U15 ( .A1(cMV1_in[6]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_h_1_n61) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_1_U14 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_1_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_1_n61), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_1_n39) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_1_U13 ( .A1(cMV1_in[5]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_h_1_n62) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_1_U12 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_1_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_1_n62), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_1_n40) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_1_U11 ( .A1(cMV1_in[4]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_h_1_n63) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_1_U10 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_1_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_1_n63), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_1_n41) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_1_U9 ( .A1(cMV1_in[3]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_h_1_n64) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_1_U8 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_1_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_1_n64), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_1_n42) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_1_U7 ( .A1(cMV1_in[2]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_h_1_n65) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_1_U6 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_1_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_1_n65), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_1_n43) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_1_U5 ( .A1(cMV1_in[1]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_h_1_n66) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_1_U4 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_1_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_1_n66), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_1_n44) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_1_U3 ( .A1(cMV1_in[0]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers1_h_1_n67) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_1_U2 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_1_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_1_n67), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_1_n45) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_1_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_1_n45), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_1__0_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_1_n56) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_1_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_1_n44), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_1__1_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_1_n55) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_1_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_1_n43), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_1__2_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_1_n54) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_1_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_1_n42), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_1__3_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_1_n53) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_1_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_1_n41), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_1__4_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_1_n52) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_1_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_1_n40), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_1__5_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_1_n51) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_1_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_1_n39), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_1__6_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_1_n50) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_1_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_1_n38), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_1__7_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_1_n49) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_1_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_1_n37), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_1__8_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_1_n48) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_1_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_1_n36), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_1__9_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_1_n47) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_1_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_1_n35), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_1_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_1__10_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_1_n46) );
  INV_X1 constructing_unit_Datapath_FaS_registers1_h_2_U24 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n33) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_2_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n66) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_2_U22 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_2_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_2_n66), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n44) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_2_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n58) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_2_U20 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_2_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_2_n58), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n36) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_2_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n59) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_2_U18 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_2_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_2_n59), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n37) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_2_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n60) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_2_U16 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_2_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_2_n60), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n38) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_2_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n63) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_2_U14 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_2_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_2_n63), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n41) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_2_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n64) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_2_U12 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_2_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_2_n64), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n42) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_2_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n65) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_2_U10 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_2_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_2_n65), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n43) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_2_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n61) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_2_U8 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_2_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_2_n61), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n39) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_2_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n62) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_2_U6 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_2_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_2_n62), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n40) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_2_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n57) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_2_U4 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_2_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_2_n57), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n35) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers1_h_2_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_h_1__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n67) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers1_h_2_U2 ( .B1(
        constructing_unit_Datapath_FaS_registers1_h_2_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers1_h_2_n67), .ZN(
        constructing_unit_Datapath_FaS_registers1_h_2_n45) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_2_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_2_n45), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_2__0_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_2_n56) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_2_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_2_n44), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_2__1_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_2_n55) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_2_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_2_n43), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_2__2_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_2_n54) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_2_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_2_n42), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_2__3_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_2_n53) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_2_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_2_n41), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_2__4_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_2_n52) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_2_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_2_n40), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_2__5_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_2_n51) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_2_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_2_n39), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_2__6_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_2_n50) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_2_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_2_n38), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_2__7_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_2_n49) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_2_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_2_n37), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_2__8_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_2_n48) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_2_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_2_n36), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_2__9_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_2_n47) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers1_h_2_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_FaS_registers1_h_2_n35), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers1_h_2_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_2__10_), .QN(
        constructing_unit_Datapath_FaS_registers1_h_2_n46) );
  INV_X1 constructing_unit_Datapath_FaS_registers2_h_1_U24 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_1_n33) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_1_U23 ( .A1(cMV2_in[10]), .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_h_1_n57) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_1_U22 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_1_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_1_n57), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_1_n35) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_1_U21 ( .A1(cMV2_in[9]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_h_1_n58) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_1_U20 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_1_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_1_n58), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_1_n36) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_1_U19 ( .A1(cMV2_in[8]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_h_1_n59) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_1_U18 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_1_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_1_n59), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_1_n37) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_1_U17 ( .A1(cMV2_in[7]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_h_1_n60) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_1_U16 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_1_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_1_n60), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_1_n38) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_1_U15 ( .A1(cMV2_in[6]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_h_1_n61) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_1_U14 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_1_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_1_n61), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_1_n39) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_1_U13 ( .A1(cMV2_in[5]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_h_1_n62) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_1_U12 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_1_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_1_n62), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_1_n40) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_1_U11 ( .A1(cMV2_in[4]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_h_1_n63) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_1_U10 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_1_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_1_n63), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_1_n41) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_1_U9 ( .A1(cMV2_in[3]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_h_1_n64) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_1_U8 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_1_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_1_n64), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_1_n42) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_1_U7 ( .A1(cMV2_in[2]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_h_1_n65) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_1_U6 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_1_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_1_n65), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_1_n43) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_1_U5 ( .A1(cMV2_in[1]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_h_1_n66) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_1_U4 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_1_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_1_n66), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_1_n44) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_1_U3 ( .A1(cMV2_in[0]), 
        .A2(1'b1), .ZN(constructing_unit_Datapath_FaS_registers2_h_1_n67) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_1_U2 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_1_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_1_n67), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_1_n45) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_1_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_1_n45), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_1__0_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_1_n56) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_1_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_1_n44), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_1__1_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_1_n55) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_1_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_1_n43), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_1__2_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_1_n54) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_1_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_1_n42), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_1__3_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_1_n53) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_1_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_1_n41), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_1__4_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_1_n52) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_1_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_1_n40), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_1__5_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_1_n51) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_1_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_1_n39), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_1__6_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_1_n50) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_1_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_1_n38), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_1__7_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_1_n49) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_1_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_1_n37), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_1__8_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_1_n48) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_1_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_1_n36), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_1__9_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_1_n47) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_1_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_1_n35), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_1_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_1__10_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_1_n46) );
  INV_X1 constructing_unit_Datapath_FaS_registers2_h_2_U24 ( .A(1'b0), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n33) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_2_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n62) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_2_U22 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_2_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_2_n62), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n40) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_2_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n57) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_2_U20 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_2_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_2_n57), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n35) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_2_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n67) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_2_U18 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_2_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_2_n67), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n45) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_2_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n66) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_2_U16 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_2_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_2_n66), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n44) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_2_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n58) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_2_U14 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_2_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_2_n58), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n36) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_2_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n59) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_2_U12 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_2_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_2_n59), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n37) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_2_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n60) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_2_U10 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_2_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_2_n60), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n38) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_2_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n63) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_2_U8 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_2_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_2_n63), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n41) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_2_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n64) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_2_U6 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_2_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_2_n64), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n42) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_2_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n65) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_2_U4 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_2_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_2_n65), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n43) );
  NAND2_X1 constructing_unit_Datapath_FaS_registers2_h_2_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_h_1__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n61) );
  OAI21_X1 constructing_unit_Datapath_FaS_registers2_h_2_U2 ( .B1(
        constructing_unit_Datapath_FaS_registers2_h_2_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_FaS_registers2_h_2_n61), .ZN(
        constructing_unit_Datapath_FaS_registers2_h_2_n39) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_2_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_2_n45), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_2__0_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_2_n56) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_2_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_2_n44), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_2__1_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_2_n55) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_2_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_2_n43), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_2__2_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_2_n54) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_2_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_2_n42), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_2__3_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_2_n53) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_2_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_2_n41), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_2__4_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_2_n52) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_2_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_2_n40), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_2__5_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_2_n51) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_2_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_2_n39), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_2__6_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_2_n50) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_2_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_2_n38), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_2__7_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_2_n49) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_2_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_2_n37), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_2__8_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_2_n48) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_2_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_2_n36), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_2__9_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_2_n47) );
  DFFR_X1 constructing_unit_Datapath_FaS_registers2_h_2_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_FaS_registers2_h_2_n35), .CK(clk), .RN(
        constructing_unit_Datapath_FaS_registers2_h_2_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_2__10_), .QN(
        constructing_unit_Datapath_FaS_registers2_h_2_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_h_3_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_3_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_h_2__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_3_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_3_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_3_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_3_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_h_2__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_3_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_3_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_3_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_3_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_h_2__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_3_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_3_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_3_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_3_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_h_2__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_3_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_3_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_3_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_3_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_h_2__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_3_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_3_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_3_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_3_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_h_2__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_3_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_3_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_3_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_3_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_h_2__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_3_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_3_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_3_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_3_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_h_2__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_3_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_3_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_3_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_3_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_h_2__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_3_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_3_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_3_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_3_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_h_2__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_3_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_3_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_3_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_3_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_h_2__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_3_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_3_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_3_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_3_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_3_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_3_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_3__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_3_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_3_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_3_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_3__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_3_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_3_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_3_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_3__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_3_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_3_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_3_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_3__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_3_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_3_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_3_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_3__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_3_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_3_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_3_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_3__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_3_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_3_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_3_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_3__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_3_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_3_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_3_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_3__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_3_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_3_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_3_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_3__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_3_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_3_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_3_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_3__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_3_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_3_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_3_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_3_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_3__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_3_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_h_4_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_4_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_h_3__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_4_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_4_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_4_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_4_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_h_3__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_4_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_4_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_4_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_4_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_h_3__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_4_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_4_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_4_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_4_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_h_3__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_4_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_4_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_4_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_4_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_h_3__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_4_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_4_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_4_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_4_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_h_3__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_4_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_4_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_4_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_4_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_h_3__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_4_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_4_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_4_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_4_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_h_3__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_4_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_4_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_4_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_4_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_h_3__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_4_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_4_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_4_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_4_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_h_3__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_4_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_4_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_4_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_4_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_h_3__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_4_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_4_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_4_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_4_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_4_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_4_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_4__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_4_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_4_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_4_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_4__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_4_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_4_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_4_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_4__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_4_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_4_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_4_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_4__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_4_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_4_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_4_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_4__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_4_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_4_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_4_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_4__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_4_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_4_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_4_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_4__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_4_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_4_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_4_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_4__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_4_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_4_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_4_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_4__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_4_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_4_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_4_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_4__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_4_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_4_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_4_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_4_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_4__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_4_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_h_5_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_5_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_h_4__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_5_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_5_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_5_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_5_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_h_4__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_5_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_5_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_5_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_5_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_h_4__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_5_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_5_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_5_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_5_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_h_4__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_5_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_5_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_5_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_5_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_h_4__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_5_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_5_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_5_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_5_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_h_4__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_5_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_5_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_5_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_5_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_h_4__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_5_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_5_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_5_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_5_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_h_4__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_5_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_5_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_5_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_5_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_h_4__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_5_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_5_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_5_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_5_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_h_4__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_5_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_5_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_5_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_5_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_h_4__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_5_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_5_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_5_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_5_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_5_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_5_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_5__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_5_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_5_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_5_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_5__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_5_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_5_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_5_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_5__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_5_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_5_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_5_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_5__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_5_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_5_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_5_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_5__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_5_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_5_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_5_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_5__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_5_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_5_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_5_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_5__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_5_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_5_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_5_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_5__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_5_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_5_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_5_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_5__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_5_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_5_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_5_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_5__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_5_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_5_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_5_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_5_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_5__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_5_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_h_6_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_6_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_h_5__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_6_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_6_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_6_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_6_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_h_5__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_6_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_6_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_6_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_6_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_h_5__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_6_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_6_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_6_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_6_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_h_5__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_6_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_6_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_6_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_6_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_h_5__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_6_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_6_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_6_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_6_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_h_5__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_6_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_6_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_6_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_6_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_h_5__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_6_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_6_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_6_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_6_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_h_5__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_6_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_6_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_6_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_6_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_h_5__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_6_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_6_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_6_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_6_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_h_5__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_6_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_6_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_6_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_6_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_h_5__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_6_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_6_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_6_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_6_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_6_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_6_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_6__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_6_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_6_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_6_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_6__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_6_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_6_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_6_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_6__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_6_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_6_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_6_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_6__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_6_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_6_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_6_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_6__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_6_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_6_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_6_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_6__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_6_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_6_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_6_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_6__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_6_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_6_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_6_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_6__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_6_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_6_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_6_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_6__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_6_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_6_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_6_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_6__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_6_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_6_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_6_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_6_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_6__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_6_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_h_7_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_7_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_h_6__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_7_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_7_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_7_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_7_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_h_6__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_7_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_7_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_7_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_7_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_h_6__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_7_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_7_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_7_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_7_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_h_6__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_7_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_7_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_7_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_7_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_h_6__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_7_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_7_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_7_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_7_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_h_6__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_7_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_7_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_7_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_7_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_h_6__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_7_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_7_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_7_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_7_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_h_6__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_7_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_7_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_7_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_7_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_h_6__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_7_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_7_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_7_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_7_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_h_6__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_7_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_7_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_7_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_7_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_h_6__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_7_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_7_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_7_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_7_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_7_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_7_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[0]), .QN(
        constructing_unit_Datapath_Middle_registers0_h_7_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_7_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_7_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[1]), .QN(
        constructing_unit_Datapath_Middle_registers0_h_7_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_7_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_7_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[2]), .QN(
        constructing_unit_Datapath_Middle_registers0_h_7_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_7_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_7_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[3]), .QN(
        constructing_unit_Datapath_Middle_registers0_h_7_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_7_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_7_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[4]), .QN(
        constructing_unit_Datapath_Middle_registers0_h_7_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_7_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_7_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[5]), .QN(
        constructing_unit_Datapath_Middle_registers0_h_7_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_7_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_7_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[6]), .QN(
        constructing_unit_Datapath_Middle_registers0_h_7_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_7_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_7_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[7]), .QN(
        constructing_unit_Datapath_Middle_registers0_h_7_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_7_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_7_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[8]), .QN(
        constructing_unit_Datapath_Middle_registers0_h_7_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_7_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_7_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[9]), .QN(
        constructing_unit_Datapath_Middle_registers0_h_7_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_7_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_7_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_7_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_ext[10]), .QN(
        constructing_unit_Datapath_Middle_registers0_h_7_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_h_8_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_8_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_h_ext[9]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_8_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_8_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_8_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_8_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_h_ext[8]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_8_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_8_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_8_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_8_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_h_ext[7]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_8_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_8_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_8_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_8_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_h_ext[6]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_8_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_8_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_8_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_8_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_h_ext[5]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_8_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_8_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_8_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_8_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_h_ext[4]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_8_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_8_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_8_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_8_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_h_ext[3]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_8_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_8_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_8_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_8_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_h_ext[2]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_8_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_8_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_8_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_8_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_h_ext[1]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_8_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_8_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_8_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_8_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_h_ext[0]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_8_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_8_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_8_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n45) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_8_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_h_ext[10]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_8_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_8_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_8_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_8_n35) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_8_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_8_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_8__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_8_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_8_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_8_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_8__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_8_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_8_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_8_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_8__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_8_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_8_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_8_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_8__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_8_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_8_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_8_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_8__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_8_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_8_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_8_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_8__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_8_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_8_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_8_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_8__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_8_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_8_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_8_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_8__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_8_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_8_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_8_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_8__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_8_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_8_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_8_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_8__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_8_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_8_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_8_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_8_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_8__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_8_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_h_9_U24 ( .A(
        constructing_unit_Datapath_n20), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_9_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_h_8__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_9_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_9_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_9_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_9_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_h_8__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_9_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_9_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_9_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_9_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_h_8__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_9_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_9_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_9_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_9_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_h_8__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_9_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_9_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_9_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_9_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_h_8__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_9_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_9_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_9_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_9_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_h_8__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_9_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_9_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_9_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_9_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_h_8__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_9_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_9_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_9_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_9_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_h_8__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_9_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_9_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_9_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_9_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_h_8__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_9_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_9_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_9_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_9_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_h_8__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_9_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_9_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_9_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_9_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_h_8__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_9_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_9_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_9_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_9_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_9_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_9_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_9__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_9_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_9_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_9_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_9__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_9_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_9_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_9_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_9__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_9_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_9_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_9_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_9__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_9_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_9_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_9_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_9__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_9_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_9_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_9_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_9__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_9_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_9_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_9_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_9__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_9_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_9_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_9_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_9__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_9_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_9_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_9_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_9__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_9_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_9_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_9_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_9__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_9_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_9_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_9_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_9_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_9__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_9_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_h_10_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_10_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_h_9__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_10_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_10_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_10_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_10_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_h_9__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_10_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_10_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_10_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_10_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_h_9__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_10_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_10_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_10_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_10_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_h_9__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_10_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_10_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_10_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_10_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_h_9__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_10_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_10_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_10_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_10_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_h_9__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_10_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_10_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_10_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_10_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_h_9__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_10_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_10_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_10_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_10_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_h_9__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_10_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_10_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_10_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_10_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_h_9__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_10_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_10_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_10_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_10_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_h_9__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_10_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_10_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_10_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_10_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_h_9__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_10_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_10_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_10_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_10_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_10_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_10_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_10__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_10_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_10_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_10_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_10__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_10_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_10_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_10_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_10__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_10_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_10_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_10_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_10__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_10_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_10_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_10_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_10__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_10_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_10_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_10_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_10__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_10_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_10_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_10_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_10__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_10_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_10_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_10_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_10__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_10_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_10_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_10_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_10__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_10_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_10_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_10_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_10__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_10_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_10_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_10_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_10_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_10__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_10_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_h_11_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_11_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_h_10__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_11_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_11_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_11_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_11_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_h_10__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_11_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_11_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_11_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_11_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_h_10__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_11_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_11_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_11_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_11_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_h_10__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_11_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_11_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_11_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_11_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_h_10__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_11_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_11_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_11_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_11_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_h_10__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_11_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_11_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_11_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_11_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_h_10__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_11_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_11_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_11_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_11_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_h_10__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_11_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_11_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_11_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_11_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_h_10__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_11_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_11_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_11_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_11_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_h_10__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_11_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_11_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_11_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_11_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_h_10__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_11_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_11_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_11_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_11_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_11_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_11_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_11__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_11_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_11_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_11_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_11__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_11_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_11_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_11_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_11__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_11_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_11_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_11_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_11__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_11_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_11_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_11_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_11__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_11_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_11_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_11_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_11__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_11_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_11_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_11_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_11__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_11_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_11_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_11_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_11__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_11_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_11_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_11_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_11__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_11_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_11_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_11_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_11__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_11_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_11_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_11_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_11_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_11__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_11_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_h_12_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_12_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_h_11__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_12_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_12_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_12_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_12_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_h_11__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_12_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_12_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_12_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_12_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_h_11__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_12_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_12_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_12_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_12_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_h_11__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_12_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_12_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_12_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_12_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_h_11__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_12_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_12_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_12_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_12_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_h_11__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_12_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_12_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_12_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_12_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_h_11__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_12_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_12_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_12_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_12_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_h_11__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_12_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_12_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_12_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_12_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_h_11__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_12_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_12_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_12_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_12_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_h_11__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_12_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_12_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_12_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_12_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_h_11__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_12_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_12_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_12_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_12_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_12_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_12_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_12__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_12_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_12_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_12_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_12__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_12_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_12_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_12_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_12__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_12_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_12_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_12_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_12__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_12_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_12_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_12_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_12__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_12_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_12_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_12_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_12__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_12_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_12_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_12_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_12__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_12_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_12_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_12_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_12__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_12_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_12_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_12_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_12__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_12_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_12_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_12_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_12__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_12_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_12_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_12_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_12_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_12__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_12_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers0_h_13_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_13_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_h_12__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_13_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_13_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_13_n57), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_13_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_h_12__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_13_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_13_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_13_n58), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_13_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_h_12__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_13_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_13_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_13_n59), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_13_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_h_12__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_13_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_13_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_13_n60), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_13_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_h_12__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_13_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_13_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_13_n61), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_13_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_h_12__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_13_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_13_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_13_n62), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_13_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_h_12__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_13_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_13_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_13_n63), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_13_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_h_12__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_13_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_13_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_13_n64), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_13_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_h_12__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_13_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_13_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_13_n65), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_13_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_h_12__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_13_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_13_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_13_n66), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers0_h_13_U3 ( .A1(
        constructing_unit_Datapath_MV0_int_h_12__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers0_h_13_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers0_h_13_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers0_h_13_n67), .ZN(
        constructing_unit_Datapath_Middle_registers0_h_13_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_13_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_13_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_13__0_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_13_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_13_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_13_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_13__1_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_13_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_13_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_13_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_13__2_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_13_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_13_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_13_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_13__3_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_13_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_13_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_13_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_13__4_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_13_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_13_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_13_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_13__5_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_13_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_13_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_13_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_13__6_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_13_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_13_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_13_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_13__7_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_13_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_13_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_13_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_13__8_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_13_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_13_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_13_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_13__9_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_13_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers0_h_13_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers0_h_13_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers0_h_13_n33), .Q(
        constructing_unit_Datapath_MV0_int_h_13__10_), .QN(
        constructing_unit_Datapath_Middle_registers0_h_13_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_3_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_3_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_h_2__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_3_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_3_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_3_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_3_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_h_2__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_3_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_3_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_3_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_3_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_h_2__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_3_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_3_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_3_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_3_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_h_2__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_3_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_3_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_3_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_3_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_h_2__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_3_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_3_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_3_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_3_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_h_2__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_3_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_3_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_3_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_3_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_h_2__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_3_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_3_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_3_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_3_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_h_2__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_3_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_3_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_3_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_3_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_h_2__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_3_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_3_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_3_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_3_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_h_2__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_3_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_3_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_3_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_3_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_h_2__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_3_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_3_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_3_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_3_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_3_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_3_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_3__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_3_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_3_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_3_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_3__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_3_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_3_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_3_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_3__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_3_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_3_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_3_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_3__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_3_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_3_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_3_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_3__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_3_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_3_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_3_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_3__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_3_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_3_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_3_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_3__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_3_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_3_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_3_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_3__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_3_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_3_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_3_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_3__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_3_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_3_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_3_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_3__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_3_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_3_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_3_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_3_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_3__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_3_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_4_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_4_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_h_3__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_4_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_4_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_4_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_4_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_h_3__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_4_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_4_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_4_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_4_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_h_3__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_4_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_4_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_4_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_4_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_h_3__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_4_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_4_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_4_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_4_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_h_3__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_4_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_4_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_4_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_4_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_h_3__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_4_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_4_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_4_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_4_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_h_3__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_4_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_4_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_4_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_4_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_h_3__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_4_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_4_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_4_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_4_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_h_3__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_4_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_4_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_4_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_4_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_h_3__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_4_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_4_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_4_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_4_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_h_3__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_4_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_4_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_4_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_4_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_4_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_4_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_4__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_4_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_4_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_4_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_4__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_4_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_4_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_4_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_4__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_4_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_4_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_4_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_4__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_4_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_4_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_4_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_4__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_4_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_4_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_4_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_4__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_4_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_4_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_4_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_4__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_4_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_4_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_4_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_4__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_4_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_4_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_4_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_4__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_4_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_4_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_4_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_4__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_4_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_4_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_4_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_4_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_4__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_4_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_5_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_5_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_h_4__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_5_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_5_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_5_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_5_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_h_4__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_5_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_5_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_5_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_5_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_h_4__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_5_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_5_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_5_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_5_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_h_4__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_5_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_5_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_5_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_5_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_h_4__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_5_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_5_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_5_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_5_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_h_4__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_5_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_5_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_5_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_5_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_h_4__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_5_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_5_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_5_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_5_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_h_4__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_5_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_5_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_5_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_5_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_h_4__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_5_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_5_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_5_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_5_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_h_4__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_5_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_5_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_5_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_5_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_h_4__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_5_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_5_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_5_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_5_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_5_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_5_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_5__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_5_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_5_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_5_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_5__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_5_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_5_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_5_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_5__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_5_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_5_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_5_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_5__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_5_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_5_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_5_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_5__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_5_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_5_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_5_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_5__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_5_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_5_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_5_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_5__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_5_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_5_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_5_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_5__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_5_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_5_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_5_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_5__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_5_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_5_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_5_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_5__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_5_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_5_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_5_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_5_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_5__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_5_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_6_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_6_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_h_5__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_6_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_6_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_6_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_6_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_h_5__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_6_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_6_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_6_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_6_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_h_5__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_6_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_6_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_6_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_6_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_h_5__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_6_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_6_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_6_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_6_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_h_5__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_6_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_6_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_6_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_6_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_h_5__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_6_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_6_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_6_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_6_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_h_5__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_6_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_6_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_6_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_6_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_h_5__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_6_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_6_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_6_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_6_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_h_5__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_6_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_6_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_6_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_6_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_h_5__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_6_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_6_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_6_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_6_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_h_5__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_6_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_6_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_6_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_6_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_6_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_6_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_6__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_6_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_6_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_6_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_6__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_6_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_6_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_6_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_6__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_6_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_6_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_6_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_6__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_6_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_6_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_6_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_6__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_6_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_6_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_6_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_6__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_6_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_6_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_6_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_6__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_6_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_6_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_6_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_6__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_6_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_6_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_6_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_6__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_6_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_6_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_6_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_6__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_6_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_6_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_6_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_6_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_6__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_6_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_7_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_7_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_h_6__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_7_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_7_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_7_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_7_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_h_6__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_7_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_7_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_7_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_7_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_h_6__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_7_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_7_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_7_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_7_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_h_6__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_7_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_7_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_7_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_7_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_h_6__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_7_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_7_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_7_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_7_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_h_6__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_7_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_7_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_7_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_7_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_h_6__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_7_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_7_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_7_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_7_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_h_6__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_7_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_7_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_7_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_7_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_h_6__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_7_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_7_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_7_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_7_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_h_6__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_7_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_7_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_7_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_7_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_h_6__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_7_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_7_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_7_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_7_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_7_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_7_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_7__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_7_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_7_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_7_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_7__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_7_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_7_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_7_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_7__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_7_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_7_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_7_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_7__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_7_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_7_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_7_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_7__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_7_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_7_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_7_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_7__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_7_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_7_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_7_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_7__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_7_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_7_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_7_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_7__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_7_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_7_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_7_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_7__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_7_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_7_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_7_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_7__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_7_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_7_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_7_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_7_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_7__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_7_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_8_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_8_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_h_7__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_8_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_8_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_8_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_8_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_h_7__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_8_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_8_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_8_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_8_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_h_7__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_8_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_8_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_8_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_8_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_h_7__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_8_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_8_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_8_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_8_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_h_7__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_8_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_8_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_8_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_8_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_h_7__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_8_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_8_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_8_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_8_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_h_7__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_8_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_8_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_8_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_8_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_h_7__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_8_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_8_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_8_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_8_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_h_7__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_8_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_8_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_8_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_8_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_h_7__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_8_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_8_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_8_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_8_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_h_7__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_8_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_8_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_8_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_8_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_8_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_8_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_8__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_8_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_8_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_8_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_8__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_8_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_8_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_8_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_8__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_8_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_8_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_8_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_8__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_8_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_8_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_8_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_8__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_8_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_8_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_8_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_8__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_8_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_8_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_8_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_8__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_8_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_8_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_8_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_8__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_8_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_8_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_8_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_8__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_8_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_8_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_8_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_8__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_8_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_8_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_8_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_8_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_8__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_8_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_9_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_9_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_h_8__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_9_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_9_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_9_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_9_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_h_8__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_9_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_9_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_9_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_9_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_h_8__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_9_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_9_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_9_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_9_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_h_8__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_9_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_9_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_9_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_9_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_h_8__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_9_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_9_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_9_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_9_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_h_8__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_9_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_9_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_9_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_9_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_h_8__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_9_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_9_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_9_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_9_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_h_8__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_9_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_9_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_9_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_9_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_h_8__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_9_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_9_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_9_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_9_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_h_8__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_9_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_9_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_9_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_9_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_h_8__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_9_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_9_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_9_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_9_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_9_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_9_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_9__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_9_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_9_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_9_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_9__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_9_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_9_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_9_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_9__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_9_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_9_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_9_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_9__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_9_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_9_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_9_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_9__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_9_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_9_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_9_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_9__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_9_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_9_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_9_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_9__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_9_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_9_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_9_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_9__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_9_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_9_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_9_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_9__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_9_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_9_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_9_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_9__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_9_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_9_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_9_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers1_9_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_9__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_9_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_10_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_10_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_h_9__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_10_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_10_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_10_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_10_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_h_9__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_10_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_10_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_10_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_10_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_h_9__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_10_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_10_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_10_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_10_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_h_9__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_10_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_10_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_10_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_10_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_h_9__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_10_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_10_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_10_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_10_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_h_9__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_10_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_10_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_10_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_10_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_h_9__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_10_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_10_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_10_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_10_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_h_9__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_10_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_10_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_10_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_10_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_h_9__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_10_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_10_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_10_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_10_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_h_9__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_10_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_10_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_10_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_10_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_h_9__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_10_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_10_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_10_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_10_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_10_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_10_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_10__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_10_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_10_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_10_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_10__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_10_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_10_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_10_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_10__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_10_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_10_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_10_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_10__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_10_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_10_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_10_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_10__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_10_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_10_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_10_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_10__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_10_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_10_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_10_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_10__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_10_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_10_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_10_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_10__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_10_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_10_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_10_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_10__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_10_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_10_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_10_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_10__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_10_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_10_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_10_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_10_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_10__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_10_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_11_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_11_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_h_10__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_11_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_11_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_11_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_11_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_h_10__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_11_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_11_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_11_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_11_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_h_10__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_11_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_11_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_11_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_11_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_h_10__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_11_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_11_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_11_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_11_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_h_10__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_11_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_11_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_11_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_11_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_h_10__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_11_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_11_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_11_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_11_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_h_10__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_11_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_11_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_11_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_11_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_h_10__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_11_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_11_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_11_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_11_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_h_10__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_11_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_11_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_11_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_11_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_h_10__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_11_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_11_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_11_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_11_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_h_10__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_11_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_11_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_11_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_11_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_11_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_11_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_11__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_11_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_11_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_11_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_11__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_11_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_11_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_11_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_11__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_11_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_11_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_11_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_11__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_11_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_11_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_11_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_11__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_11_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_11_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_11_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_11__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_11_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_11_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_11_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_11__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_11_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_11_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_11_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_11__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_11_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_11_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_11_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_11__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_11_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_11_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_11_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_11__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_11_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_11_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_11_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_11_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_11__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_11_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_12_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_12_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_h_11__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_12_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_12_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_12_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_12_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_h_11__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_12_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_12_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_12_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_12_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_h_11__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_12_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_12_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_12_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_12_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_h_11__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_12_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_12_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_12_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_12_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_h_11__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_12_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_12_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_12_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_12_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_h_11__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_12_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_12_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_12_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_12_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_h_11__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_12_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_12_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_12_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_12_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_h_11__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_12_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_12_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_12_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_12_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_h_11__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_12_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_12_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_12_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_12_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_h_11__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_12_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_12_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_12_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_12_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_h_11__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_12_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_12_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_12_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_12_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_12_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_12_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_12__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_12_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_12_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_12_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_12__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_12_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_12_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_12_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_12__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_12_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_12_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_12_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_12__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_12_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_12_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_12_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_12__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_12_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_12_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_12_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_12__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_12_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_12_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_12_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_12__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_12_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_12_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_12_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_12__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_12_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_12_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_12_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_12__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_12_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_12_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_12_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_12__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_12_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_12_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_12_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_12_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_12__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_12_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers1_13_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_13_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_h_12__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_13_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers1_13_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_13_n57), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_13_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_h_12__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_13_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers1_13_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_13_n58), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_13_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_h_12__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_13_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers1_13_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_13_n59), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_13_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_h_12__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_13_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers1_13_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_13_n60), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_13_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_h_12__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_13_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers1_13_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_13_n61), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_13_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_h_12__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_13_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers1_13_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_13_n62), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_13_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_h_12__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_13_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers1_13_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_13_n63), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_13_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_h_12__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_13_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers1_13_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_13_n64), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_13_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_h_12__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_13_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers1_13_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_13_n65), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_13_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_h_12__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_13_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers1_13_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_13_n66), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers1_13_U3 ( .A1(
        constructing_unit_Datapath_MV1_int_h_12__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers1_13_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers1_13_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers1_13_n67), .ZN(
        constructing_unit_Datapath_Middle_registers1_13_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_13_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_13_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_13__0_), .QN(
        constructing_unit_Datapath_Middle_registers1_13_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_13_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_13_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_13__1_), .QN(
        constructing_unit_Datapath_Middle_registers1_13_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_13_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_13_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_13__2_), .QN(
        constructing_unit_Datapath_Middle_registers1_13_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_13_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_13_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_13__3_), .QN(
        constructing_unit_Datapath_Middle_registers1_13_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_13_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_13_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_13__4_), .QN(
        constructing_unit_Datapath_Middle_registers1_13_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_13_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_13_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_13__5_), .QN(
        constructing_unit_Datapath_Middle_registers1_13_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_13_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_13_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_13__6_), .QN(
        constructing_unit_Datapath_Middle_registers1_13_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_13_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_13_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_13__7_), .QN(
        constructing_unit_Datapath_Middle_registers1_13_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_13_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_13_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_13__8_), .QN(
        constructing_unit_Datapath_Middle_registers1_13_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_13_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_13_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_13__9_), .QN(
        constructing_unit_Datapath_Middle_registers1_13_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers1_13_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers1_13_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers1_13_n33), .Q(
        constructing_unit_Datapath_MV1_int_h_13__10_), .QN(
        constructing_unit_Datapath_Middle_registers1_13_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_3_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_3_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_h_2__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_3_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_3_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_3_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_3_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_h_2__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_3_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_3_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_3_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_3_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_h_2__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_3_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_3_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_3_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_3_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_h_2__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_3_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_3_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_3_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_3_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_h_2__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_3_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_3_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_3_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_3_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_h_2__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_3_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_3_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_3_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_3_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_h_2__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_3_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_3_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_3_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_3_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_h_2__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_3_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_3_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_3_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_3_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_h_2__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_3_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_3_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_3_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_3_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_h_2__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_3_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_3_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_3_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_3_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_h_2__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_3_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_3_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_3_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_3_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_3_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_3_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_3__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_3_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_3_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_3_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_3__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_3_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_3_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_3_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_3__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_3_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_3_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_3_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_3__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_3_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_3_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_3_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_3__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_3_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_3_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_3_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_3__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_3_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_3_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_3_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_3__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_3_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_3_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_3_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_3__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_3_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_3_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_3_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_3__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_3_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_3_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_3_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_3__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_3_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_3_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_3_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_3_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_3__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_3_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_4_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_4_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_h_3__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_4_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_4_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_4_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_4_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_h_3__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_4_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_4_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_4_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_4_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_h_3__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_4_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_4_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_4_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_4_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_h_3__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_4_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_4_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_4_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_4_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_h_3__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_4_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_4_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_4_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_4_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_h_3__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_4_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_4_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_4_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_4_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_h_3__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_4_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_4_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_4_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_4_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_h_3__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_4_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_4_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_4_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_4_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_h_3__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_4_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_4_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_4_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_4_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_h_3__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_4_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_4_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_4_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_4_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_h_3__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_4_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_4_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_4_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_4_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_4_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_4_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_4__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_4_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_4_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_4_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_4__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_4_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_4_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_4_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_4__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_4_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_4_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_4_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_4__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_4_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_4_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_4_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_4__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_4_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_4_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_4_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_4__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_4_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_4_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_4_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_4__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_4_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_4_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_4_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_4__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_4_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_4_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_4_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_4__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_4_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_4_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_4_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_4__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_4_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_4_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_4_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_4_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_4__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_4_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_5_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_5_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_h_4__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_5_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_5_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_5_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_5_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_h_4__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_5_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_5_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_5_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_5_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_h_4__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_5_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_5_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_5_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_5_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_h_4__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_5_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_5_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_5_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_5_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_h_4__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_5_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_5_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_5_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_5_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_h_4__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_5_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_5_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_5_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_5_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_h_4__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_5_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_5_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_5_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_5_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_h_4__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_5_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_5_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_5_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_5_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_h_4__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_5_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_5_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_5_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_5_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_h_4__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_5_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_5_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_5_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_5_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_h_4__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_5_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_5_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_5_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_5_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_5_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_5_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_5__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_5_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_5_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_5_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_5__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_5_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_5_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_5_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_5__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_5_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_5_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_5_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_5__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_5_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_5_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_5_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_5__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_5_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_5_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_5_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_5__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_5_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_5_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_5_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_5__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_5_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_5_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_5_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_5__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_5_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_5_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_5_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_5__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_5_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_5_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_5_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_5__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_5_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_5_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_5_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_5_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_5__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_5_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_6_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_6_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_h_5__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_6_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_6_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_6_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_6_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_h_5__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_6_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_6_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_6_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_6_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_h_5__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_6_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_6_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_6_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_6_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_h_5__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_6_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_6_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_6_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_6_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_h_5__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_6_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_6_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_6_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_6_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_h_5__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_6_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_6_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_6_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_6_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_h_5__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_6_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_6_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_6_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_6_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_h_5__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_6_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_6_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_6_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_6_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_h_5__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_6_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_6_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_6_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_6_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_h_5__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_6_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_6_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_6_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_6_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_h_5__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_6_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_6_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_6_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_6_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_6_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_6_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_6__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_6_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_6_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_6_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_6__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_6_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_6_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_6_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_6__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_6_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_6_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_6_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_6__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_6_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_6_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_6_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_6__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_6_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_6_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_6_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_6__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_6_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_6_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_6_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_6__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_6_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_6_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_6_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_6__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_6_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_6_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_6_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_6__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_6_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_6_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_6_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_6__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_6_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_6_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_6_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_6_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_6__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_6_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_7_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_7_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_h_6__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_7_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_7_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_7_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_7_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_h_6__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_7_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_7_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_7_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_7_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_h_6__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_7_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_7_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_7_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_7_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_h_6__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_7_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_7_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_7_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_7_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_h_6__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_7_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_7_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_7_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_7_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_h_6__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_7_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_7_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_7_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_7_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_h_6__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_7_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_7_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_7_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_7_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_h_6__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_7_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_7_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_7_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_7_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_h_6__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_7_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_7_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_7_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_7_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_h_6__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_7_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_7_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_7_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_7_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_h_6__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_7_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_7_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_7_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_7_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_7_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_7_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_7__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_7_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_7_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_7_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_7__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_7_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_7_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_7_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_7__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_7_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_7_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_7_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_7__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_7_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_7_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_7_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_7__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_7_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_7_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_7_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_7__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_7_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_7_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_7_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_7__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_7_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_7_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_7_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_7__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_7_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_7_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_7_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_7__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_7_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_7_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_7_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_7__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_7_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_7_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_7_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_7_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_7__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_7_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_8_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_8_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_h_7__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_8_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_8_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_8_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_8_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_h_7__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_8_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_8_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_8_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_8_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_h_7__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_8_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_8_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_8_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_8_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_h_7__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_8_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_8_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_8_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_8_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_h_7__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_8_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_8_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_8_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_8_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_h_7__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_8_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_8_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_8_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_8_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_h_7__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_8_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_8_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_8_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_8_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_h_7__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_8_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_8_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_8_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_8_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_h_7__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_8_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_8_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_8_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_8_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_h_7__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_8_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_8_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_8_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_8_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_h_7__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_8_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_8_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_8_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_8_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_8_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_8_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[0]), .QN(
        constructing_unit_Datapath_Middle_registers2_8_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_8_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_8_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[1]), .QN(
        constructing_unit_Datapath_Middle_registers2_8_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_8_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_8_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[2]), .QN(
        constructing_unit_Datapath_Middle_registers2_8_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_8_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_8_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[3]), .QN(
        constructing_unit_Datapath_Middle_registers2_8_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_8_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_8_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[4]), .QN(
        constructing_unit_Datapath_Middle_registers2_8_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_8_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_8_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[5]), .QN(
        constructing_unit_Datapath_Middle_registers2_8_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_8_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_8_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[6]), .QN(
        constructing_unit_Datapath_Middle_registers2_8_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_8_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_8_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[7]), .QN(
        constructing_unit_Datapath_Middle_registers2_8_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_8_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_8_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[8]), .QN(
        constructing_unit_Datapath_Middle_registers2_8_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_8_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_8_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[9]), .QN(
        constructing_unit_Datapath_Middle_registers2_8_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_8_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_8_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_8_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_ext[10]), .QN(
        constructing_unit_Datapath_Middle_registers2_8_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_9_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_9_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_h_ext[9]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_9_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_9_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_9_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_9_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_h_ext[8]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_9_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_9_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_9_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_9_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_h_ext[7]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_9_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_9_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_9_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_9_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_h_ext[6]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_9_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_9_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_9_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_9_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_h_ext[5]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_9_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_9_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_9_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_9_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_h_ext[4]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_9_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_9_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_9_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_9_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_h_ext[3]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_9_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_9_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_9_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_9_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_h_ext[2]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_9_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_9_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_9_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_9_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_h_ext[1]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_9_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_9_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_9_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_9_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_h_ext[0]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_9_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_9_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_9_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n45) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_9_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_h_ext[10]), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_9_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_9_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_9_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_9_n35) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_9_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_9_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_9__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_9_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_9_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_9_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_9__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_9_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_9_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_9_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_9__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_9_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_9_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_9_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_9__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_9_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_9_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_9_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_9__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_9_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_9_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_9_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_9__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_9_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_9_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_9_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_9__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_9_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_9_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_9_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_9__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_9_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_9_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_9_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_9__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_9_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_9_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_9_n36), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_9__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_9_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_9_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_9_n35), .CK(clk), .RN(
        constructing_unit_Datapath_Middle_registers2_9_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_9__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_9_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_10_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_10_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_h_9__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_10_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_10_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_10_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_10_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_h_9__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_10_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_10_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_10_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_10_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_h_9__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_10_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_10_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_10_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_10_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_h_9__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_10_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_10_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_10_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_10_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_h_9__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_10_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_10_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_10_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_10_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_h_9__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_10_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_10_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_10_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_10_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_h_9__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_10_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_10_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_10_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_10_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_h_9__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_10_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_10_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_10_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_10_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_h_9__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_10_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_10_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_10_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_10_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_h_9__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_10_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_10_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_10_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_10_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_h_9__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_10_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_10_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_10_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_10_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_10_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_10_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_10__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_10_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_10_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_10_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_10__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_10_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_10_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_10_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_10__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_10_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_10_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_10_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_10__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_10_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_10_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_10_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_10__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_10_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_10_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_10_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_10__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_10_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_10_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_10_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_10__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_10_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_10_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_10_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_10__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_10_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_10_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_10_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_10__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_10_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_10_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_10_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_10__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_10_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_10_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_10_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_10_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_10__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_10_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_11_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_11_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_h_10__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_11_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_11_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_11_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_11_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_h_10__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_11_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_11_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_11_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_11_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_h_10__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_11_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_11_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_11_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_11_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_h_10__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_11_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_11_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_11_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_11_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_h_10__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_11_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_11_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_11_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_11_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_h_10__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_11_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_11_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_11_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_11_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_h_10__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_11_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_11_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_11_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_11_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_h_10__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_11_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_11_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_11_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_11_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_h_10__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_11_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_11_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_11_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_11_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_h_10__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_11_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_11_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_11_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_11_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_h_10__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_11_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_11_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_11_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_11_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_11_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_11_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_11__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_11_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_11_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_11_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_11__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_11_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_11_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_11_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_11__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_11_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_11_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_11_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_11__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_11_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_11_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_11_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_11__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_11_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_11_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_11_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_11__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_11_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_11_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_11_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_11__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_11_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_11_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_11_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_11__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_11_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_11_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_11_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_11__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_11_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_11_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_11_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_11__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_11_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_11_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_11_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_11_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_11__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_11_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_12_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_12_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_h_11__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_12_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_12_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_12_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_12_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_h_11__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_12_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_12_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_12_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_12_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_h_11__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_12_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_12_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_12_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_12_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_h_11__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_12_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_12_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_12_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_12_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_h_11__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_12_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_12_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_12_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_12_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_h_11__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_12_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_12_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_12_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_12_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_h_11__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_12_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_12_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_12_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_12_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_h_11__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_12_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_12_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_12_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_12_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_h_11__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_12_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_12_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_12_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_12_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_h_11__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_12_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_12_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_12_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_12_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_h_11__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_12_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_12_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_12_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_12_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_12_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_12_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_12__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_12_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_12_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_12_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_12__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_12_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_12_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_12_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_12__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_12_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_12_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_12_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_12__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_12_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_12_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_12_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_12__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_12_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_12_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_12_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_12__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_12_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_12_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_12_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_12__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_12_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_12_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_12_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_12__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_12_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_12_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_12_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_12__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_12_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_12_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_12_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_12__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_12_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_12_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_12_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_12_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_12__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_12_n46) );
  INV_X1 constructing_unit_Datapath_Middle_registers2_13_U24 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n33) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_13_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_h_12__10_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n57) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_13_U22 ( .B1(
        constructing_unit_Datapath_Middle_registers2_13_n46), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_13_n57), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n35) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_13_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_h_12__9_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n58) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_13_U20 ( .B1(
        constructing_unit_Datapath_Middle_registers2_13_n47), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_13_n58), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n36) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_13_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_h_12__8_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n59) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_13_U18 ( .B1(
        constructing_unit_Datapath_Middle_registers2_13_n48), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_13_n59), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n37) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_13_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_h_12__7_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n60) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_13_U16 ( .B1(
        constructing_unit_Datapath_Middle_registers2_13_n49), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_13_n60), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n38) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_13_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_h_12__6_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n61) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_13_U14 ( .B1(
        constructing_unit_Datapath_Middle_registers2_13_n50), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_13_n61), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n39) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_13_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_h_12__5_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n62) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_13_U12 ( .B1(
        constructing_unit_Datapath_Middle_registers2_13_n51), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_13_n62), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n40) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_13_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_h_12__4_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n63) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_13_U10 ( .B1(
        constructing_unit_Datapath_Middle_registers2_13_n52), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_13_n63), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n41) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_13_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_h_12__3_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n64) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_13_U8 ( .B1(
        constructing_unit_Datapath_Middle_registers2_13_n53), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_13_n64), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n42) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_13_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_h_12__2_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n65) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_13_U6 ( .B1(
        constructing_unit_Datapath_Middle_registers2_13_n54), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_13_n65), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n43) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_13_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_h_12__1_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n66) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_13_U4 ( .B1(
        constructing_unit_Datapath_Middle_registers2_13_n55), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_13_n66), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n44) );
  NAND2_X1 constructing_unit_Datapath_Middle_registers2_13_U3 ( .A1(
        constructing_unit_Datapath_MV2_int_h_12__0_), .A2(1'b1), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n67) );
  OAI21_X1 constructing_unit_Datapath_Middle_registers2_13_U2 ( .B1(
        constructing_unit_Datapath_Middle_registers2_13_n56), .B2(1'b1), .A(
        constructing_unit_Datapath_Middle_registers2_13_n67), .ZN(
        constructing_unit_Datapath_Middle_registers2_13_n45) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_13_MV_out_int_reg_0_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_13_n45), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_13__0_), .QN(
        constructing_unit_Datapath_Middle_registers2_13_n56) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_13_MV_out_int_reg_1_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_13_n44), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_13__1_), .QN(
        constructing_unit_Datapath_Middle_registers2_13_n55) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_13_MV_out_int_reg_2_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_13_n43), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_13__2_), .QN(
        constructing_unit_Datapath_Middle_registers2_13_n54) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_13_MV_out_int_reg_3_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_13_n42), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_13__3_), .QN(
        constructing_unit_Datapath_Middle_registers2_13_n53) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_13_MV_out_int_reg_4_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_13_n41), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_13__4_), .QN(
        constructing_unit_Datapath_Middle_registers2_13_n52) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_13_MV_out_int_reg_5_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_13_n40), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_13__5_), .QN(
        constructing_unit_Datapath_Middle_registers2_13_n51) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_13_MV_out_int_reg_6_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_13_n39), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_13__6_), .QN(
        constructing_unit_Datapath_Middle_registers2_13_n50) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_13_MV_out_int_reg_7_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_13_n38), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_13__7_), .QN(
        constructing_unit_Datapath_Middle_registers2_13_n49) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_13_MV_out_int_reg_8_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_13_n37), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_13__8_), .QN(
        constructing_unit_Datapath_Middle_registers2_13_n48) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_13_MV_out_int_reg_9_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_13_n36), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_13__9_), .QN(
        constructing_unit_Datapath_Middle_registers2_13_n47) );
  DFFR_X1 constructing_unit_Datapath_Middle_registers2_13_MV_out_int_reg_10_ ( 
        .D(constructing_unit_Datapath_Middle_registers2_13_n35), .CK(clk), 
        .RN(constructing_unit_Datapath_Middle_registers2_13_n33), .Q(
        constructing_unit_Datapath_MV2_int_h_13__10_), .QN(
        constructing_unit_Datapath_Middle_registers2_13_n46) );
  INV_X1 constructing_unit_Datapath_Last_register0_h_U26 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Last_register0_h_n36) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_h_U25 ( .A1(
        constructing_unit_Datapath_MV0_int_h_13__9_), .A2(
        constructing_unit_Datapath_Last_register0_h_n33), .ZN(
        constructing_unit_Datapath_Last_register0_h_n60) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_h_U24 ( .B1(
        constructing_unit_Datapath_Last_register0_h_n49), .B2(
        constructing_unit_Datapath_Last_register0_h_n35), .A(
        constructing_unit_Datapath_Last_register0_h_n60), .ZN(
        constructing_unit_Datapath_Last_register0_h_n38) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_h_U23 ( .A1(
        constructing_unit_Datapath_MV0_int_h_13__8_), .A2(
        constructing_unit_Datapath_Last_register0_h_n33), .ZN(
        constructing_unit_Datapath_Last_register0_h_n61) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_h_U22 ( .B1(
        constructing_unit_Datapath_Last_register0_h_n50), .B2(
        constructing_unit_Datapath_Last_register0_h_n35), .A(
        constructing_unit_Datapath_Last_register0_h_n61), .ZN(
        constructing_unit_Datapath_Last_register0_h_n39) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_h_U21 ( .A1(
        constructing_unit_Datapath_MV0_int_h_13__7_), .A2(
        constructing_unit_Datapath_Last_register0_h_n33), .ZN(
        constructing_unit_Datapath_Last_register0_h_n62) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_h_U20 ( .B1(
        constructing_unit_Datapath_Last_register0_h_n51), .B2(
        constructing_unit_Datapath_Last_register0_h_n35), .A(
        constructing_unit_Datapath_Last_register0_h_n62), .ZN(
        constructing_unit_Datapath_Last_register0_h_n40) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_h_U19 ( .A1(
        constructing_unit_Datapath_MV0_int_h_13__6_), .A2(
        constructing_unit_Datapath_Last_register0_h_n33), .ZN(
        constructing_unit_Datapath_Last_register0_h_n63) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_h_U18 ( .B1(
        constructing_unit_Datapath_Last_register0_h_n52), .B2(
        constructing_unit_Datapath_Last_register0_h_n35), .A(
        constructing_unit_Datapath_Last_register0_h_n63), .ZN(
        constructing_unit_Datapath_Last_register0_h_n41) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_h_U17 ( .A1(
        constructing_unit_Datapath_MV0_int_h_13__5_), .A2(
        constructing_unit_Datapath_Last_register0_h_n33), .ZN(
        constructing_unit_Datapath_Last_register0_h_n64) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_h_U16 ( .B1(
        constructing_unit_Datapath_Last_register0_h_n53), .B2(
        constructing_unit_Datapath_Last_register0_h_n35), .A(
        constructing_unit_Datapath_Last_register0_h_n64), .ZN(
        constructing_unit_Datapath_Last_register0_h_n42) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_h_U15 ( .A1(
        constructing_unit_Datapath_MV0_int_h_13__4_), .A2(
        constructing_unit_Datapath_Last_register0_h_n33), .ZN(
        constructing_unit_Datapath_Last_register0_h_n65) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_h_U14 ( .B1(
        constructing_unit_Datapath_Last_register0_h_n54), .B2(
        constructing_unit_Datapath_Last_register0_h_n35), .A(
        constructing_unit_Datapath_Last_register0_h_n65), .ZN(
        constructing_unit_Datapath_Last_register0_h_n43) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_h_U13 ( .A1(
        constructing_unit_Datapath_MV0_int_h_13__3_), .A2(
        constructing_unit_Datapath_Last_register0_h_n33), .ZN(
        constructing_unit_Datapath_Last_register0_h_n66) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_h_U12 ( .B1(
        constructing_unit_Datapath_Last_register0_h_n55), .B2(
        constructing_unit_Datapath_Last_register0_h_n35), .A(
        constructing_unit_Datapath_Last_register0_h_n66), .ZN(
        constructing_unit_Datapath_Last_register0_h_n44) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_h_U11 ( .A1(
        constructing_unit_Datapath_MV0_int_h_13__2_), .A2(
        constructing_unit_Datapath_Last_register0_h_n33), .ZN(
        constructing_unit_Datapath_Last_register0_h_n67) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_h_U10 ( .B1(
        constructing_unit_Datapath_Last_register0_h_n56), .B2(
        constructing_unit_Datapath_Last_register0_h_n35), .A(
        constructing_unit_Datapath_Last_register0_h_n67), .ZN(
        constructing_unit_Datapath_Last_register0_h_n45) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_h_U9 ( .A1(
        constructing_unit_Datapath_MV0_int_h_13__1_), .A2(
        constructing_unit_Datapath_Last_register0_h_n33), .ZN(
        constructing_unit_Datapath_Last_register0_h_n68) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_h_U8 ( .B1(
        constructing_unit_Datapath_Last_register0_h_n57), .B2(
        constructing_unit_Datapath_Last_register0_h_n35), .A(
        constructing_unit_Datapath_Last_register0_h_n68), .ZN(
        constructing_unit_Datapath_Last_register0_h_n46) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_h_U7 ( .A1(
        constructing_unit_Datapath_MV0_int_h_13__0_), .A2(
        constructing_unit_Datapath_Last_register0_h_n33), .ZN(
        constructing_unit_Datapath_Last_register0_h_n69) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_h_U6 ( .B1(
        constructing_unit_Datapath_Last_register0_h_n58), .B2(
        constructing_unit_Datapath_Last_register0_h_n35), .A(
        constructing_unit_Datapath_Last_register0_h_n69), .ZN(
        constructing_unit_Datapath_Last_register0_h_n47) );
  NAND2_X1 constructing_unit_Datapath_Last_register0_h_U5 ( .A1(
        constructing_unit_Datapath_MV0_int_h_13__10_), .A2(
        constructing_unit_Datapath_Last_register0_h_n33), .ZN(
        constructing_unit_Datapath_Last_register0_h_n59) );
  OAI21_X1 constructing_unit_Datapath_Last_register0_h_U4 ( .B1(
        constructing_unit_Datapath_Last_register0_h_n48), .B2(
        constructing_unit_Datapath_Last_register0_h_n33), .A(
        constructing_unit_Datapath_Last_register0_h_n59), .ZN(
        constructing_unit_Datapath_Last_register0_h_n37) );
  BUF_X1 constructing_unit_Datapath_Last_register0_h_U3 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_Last_register0_h_n35) );
  BUF_X1 constructing_unit_Datapath_Last_register0_h_U2 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_Last_register0_h_n33) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_h_MV_out_int_reg_0_ ( .D(
        constructing_unit_Datapath_Last_register0_h_n47), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_h_n36), .Q(MVP0[0]), .QN(
        constructing_unit_Datapath_Last_register0_h_n58) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_h_MV_out_int_reg_1_ ( .D(
        constructing_unit_Datapath_Last_register0_h_n46), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_h_n36), .Q(MVP0[1]), .QN(
        constructing_unit_Datapath_Last_register0_h_n57) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_h_MV_out_int_reg_2_ ( .D(
        constructing_unit_Datapath_Last_register0_h_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_h_n36), .Q(MVP0[2]), .QN(
        constructing_unit_Datapath_Last_register0_h_n56) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_h_MV_out_int_reg_3_ ( .D(
        constructing_unit_Datapath_Last_register0_h_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_h_n36), .Q(MVP0[3]), .QN(
        constructing_unit_Datapath_Last_register0_h_n55) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_h_MV_out_int_reg_4_ ( .D(
        constructing_unit_Datapath_Last_register0_h_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_h_n36), .Q(MVP0[4]), .QN(
        constructing_unit_Datapath_Last_register0_h_n54) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_h_MV_out_int_reg_5_ ( .D(
        constructing_unit_Datapath_Last_register0_h_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_h_n36), .Q(MVP0[5]), .QN(
        constructing_unit_Datapath_Last_register0_h_n53) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_h_MV_out_int_reg_6_ ( .D(
        constructing_unit_Datapath_Last_register0_h_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_h_n36), .Q(MVP0[6]), .QN(
        constructing_unit_Datapath_Last_register0_h_n52) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_h_MV_out_int_reg_7_ ( .D(
        constructing_unit_Datapath_Last_register0_h_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_h_n36), .Q(MVP0[7]), .QN(
        constructing_unit_Datapath_Last_register0_h_n51) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_h_MV_out_int_reg_8_ ( .D(
        constructing_unit_Datapath_Last_register0_h_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_h_n36), .Q(MVP0[8]), .QN(
        constructing_unit_Datapath_Last_register0_h_n50) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_h_MV_out_int_reg_9_ ( .D(
        constructing_unit_Datapath_Last_register0_h_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_h_n36), .Q(MVP0[9]), .QN(
        constructing_unit_Datapath_Last_register0_h_n49) );
  DFFR_X1 constructing_unit_Datapath_Last_register0_h_MV_out_int_reg_10_ ( .D(
        constructing_unit_Datapath_Last_register0_h_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register0_h_n36), .Q(MVP0[10]), .QN(
        constructing_unit_Datapath_Last_register0_h_n48) );
  INV_X1 constructing_unit_Datapath_Last_register1_h_U26 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Last_register1_h_n36) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_h_U25 ( .A1(
        constructing_unit_Datapath_MV1_int_h_13__9_), .A2(
        constructing_unit_Datapath_Last_register1_h_n33), .ZN(
        constructing_unit_Datapath_Last_register1_h_n60) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_h_U24 ( .B1(
        constructing_unit_Datapath_Last_register1_h_n49), .B2(
        constructing_unit_Datapath_Last_register1_h_n35), .A(
        constructing_unit_Datapath_Last_register1_h_n60), .ZN(
        constructing_unit_Datapath_Last_register1_h_n38) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_h_U23 ( .A1(
        constructing_unit_Datapath_MV1_int_h_13__8_), .A2(
        constructing_unit_Datapath_Last_register1_h_n33), .ZN(
        constructing_unit_Datapath_Last_register1_h_n61) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_h_U22 ( .B1(
        constructing_unit_Datapath_Last_register1_h_n50), .B2(
        constructing_unit_Datapath_Last_register1_h_n35), .A(
        constructing_unit_Datapath_Last_register1_h_n61), .ZN(
        constructing_unit_Datapath_Last_register1_h_n39) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_h_U21 ( .A1(
        constructing_unit_Datapath_MV1_int_h_13__7_), .A2(
        constructing_unit_Datapath_Last_register1_h_n33), .ZN(
        constructing_unit_Datapath_Last_register1_h_n62) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_h_U20 ( .B1(
        constructing_unit_Datapath_Last_register1_h_n51), .B2(
        constructing_unit_Datapath_Last_register1_h_n35), .A(
        constructing_unit_Datapath_Last_register1_h_n62), .ZN(
        constructing_unit_Datapath_Last_register1_h_n40) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_h_U19 ( .A1(
        constructing_unit_Datapath_MV1_int_h_13__6_), .A2(
        constructing_unit_Datapath_Last_register1_h_n33), .ZN(
        constructing_unit_Datapath_Last_register1_h_n63) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_h_U18 ( .B1(
        constructing_unit_Datapath_Last_register1_h_n52), .B2(
        constructing_unit_Datapath_Last_register1_h_n35), .A(
        constructing_unit_Datapath_Last_register1_h_n63), .ZN(
        constructing_unit_Datapath_Last_register1_h_n41) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_h_U17 ( .A1(
        constructing_unit_Datapath_MV1_int_h_13__5_), .A2(
        constructing_unit_Datapath_Last_register1_h_n33), .ZN(
        constructing_unit_Datapath_Last_register1_h_n64) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_h_U16 ( .B1(
        constructing_unit_Datapath_Last_register1_h_n53), .B2(
        constructing_unit_Datapath_Last_register1_h_n35), .A(
        constructing_unit_Datapath_Last_register1_h_n64), .ZN(
        constructing_unit_Datapath_Last_register1_h_n42) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_h_U15 ( .A1(
        constructing_unit_Datapath_MV1_int_h_13__4_), .A2(
        constructing_unit_Datapath_Last_register1_h_n33), .ZN(
        constructing_unit_Datapath_Last_register1_h_n65) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_h_U14 ( .B1(
        constructing_unit_Datapath_Last_register1_h_n54), .B2(
        constructing_unit_Datapath_Last_register1_h_n35), .A(
        constructing_unit_Datapath_Last_register1_h_n65), .ZN(
        constructing_unit_Datapath_Last_register1_h_n43) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_h_U13 ( .A1(
        constructing_unit_Datapath_MV1_int_h_13__3_), .A2(
        constructing_unit_Datapath_Last_register1_h_n33), .ZN(
        constructing_unit_Datapath_Last_register1_h_n66) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_h_U12 ( .B1(
        constructing_unit_Datapath_Last_register1_h_n55), .B2(
        constructing_unit_Datapath_Last_register1_h_n35), .A(
        constructing_unit_Datapath_Last_register1_h_n66), .ZN(
        constructing_unit_Datapath_Last_register1_h_n44) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_h_U11 ( .A1(
        constructing_unit_Datapath_MV1_int_h_13__2_), .A2(
        constructing_unit_Datapath_Last_register1_h_n33), .ZN(
        constructing_unit_Datapath_Last_register1_h_n67) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_h_U10 ( .B1(
        constructing_unit_Datapath_Last_register1_h_n56), .B2(
        constructing_unit_Datapath_Last_register1_h_n35), .A(
        constructing_unit_Datapath_Last_register1_h_n67), .ZN(
        constructing_unit_Datapath_Last_register1_h_n45) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_h_U9 ( .A1(
        constructing_unit_Datapath_MV1_int_h_13__1_), .A2(
        constructing_unit_Datapath_Last_register1_h_n33), .ZN(
        constructing_unit_Datapath_Last_register1_h_n68) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_h_U8 ( .B1(
        constructing_unit_Datapath_Last_register1_h_n57), .B2(
        constructing_unit_Datapath_Last_register1_h_n35), .A(
        constructing_unit_Datapath_Last_register1_h_n68), .ZN(
        constructing_unit_Datapath_Last_register1_h_n46) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_h_U7 ( .A1(
        constructing_unit_Datapath_MV1_int_h_13__0_), .A2(
        constructing_unit_Datapath_Last_register1_h_n33), .ZN(
        constructing_unit_Datapath_Last_register1_h_n69) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_h_U6 ( .B1(
        constructing_unit_Datapath_Last_register1_h_n58), .B2(
        constructing_unit_Datapath_Last_register1_h_n35), .A(
        constructing_unit_Datapath_Last_register1_h_n69), .ZN(
        constructing_unit_Datapath_Last_register1_h_n47) );
  NAND2_X1 constructing_unit_Datapath_Last_register1_h_U5 ( .A1(
        constructing_unit_Datapath_MV1_int_h_13__10_), .A2(
        constructing_unit_Datapath_Last_register1_h_n33), .ZN(
        constructing_unit_Datapath_Last_register1_h_n59) );
  OAI21_X1 constructing_unit_Datapath_Last_register1_h_U4 ( .B1(
        constructing_unit_Datapath_Last_register1_h_n48), .B2(
        constructing_unit_Datapath_Last_register1_h_n33), .A(
        constructing_unit_Datapath_Last_register1_h_n59), .ZN(
        constructing_unit_Datapath_Last_register1_h_n37) );
  BUF_X1 constructing_unit_Datapath_Last_register1_h_U3 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_Last_register1_h_n35) );
  BUF_X1 constructing_unit_Datapath_Last_register1_h_U2 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_Last_register1_h_n33) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_h_MV_out_int_reg_0_ ( .D(
        constructing_unit_Datapath_Last_register1_h_n47), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_h_n36), .Q(MVP1[0]), .QN(
        constructing_unit_Datapath_Last_register1_h_n58) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_h_MV_out_int_reg_1_ ( .D(
        constructing_unit_Datapath_Last_register1_h_n46), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_h_n36), .Q(MVP1[1]), .QN(
        constructing_unit_Datapath_Last_register1_h_n57) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_h_MV_out_int_reg_2_ ( .D(
        constructing_unit_Datapath_Last_register1_h_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_h_n36), .Q(MVP1[2]), .QN(
        constructing_unit_Datapath_Last_register1_h_n56) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_h_MV_out_int_reg_3_ ( .D(
        constructing_unit_Datapath_Last_register1_h_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_h_n36), .Q(MVP1[3]), .QN(
        constructing_unit_Datapath_Last_register1_h_n55) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_h_MV_out_int_reg_4_ ( .D(
        constructing_unit_Datapath_Last_register1_h_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_h_n36), .Q(MVP1[4]), .QN(
        constructing_unit_Datapath_Last_register1_h_n54) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_h_MV_out_int_reg_5_ ( .D(
        constructing_unit_Datapath_Last_register1_h_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_h_n36), .Q(MVP1[5]), .QN(
        constructing_unit_Datapath_Last_register1_h_n53) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_h_MV_out_int_reg_6_ ( .D(
        constructing_unit_Datapath_Last_register1_h_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_h_n36), .Q(MVP1[6]), .QN(
        constructing_unit_Datapath_Last_register1_h_n52) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_h_MV_out_int_reg_7_ ( .D(
        constructing_unit_Datapath_Last_register1_h_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_h_n36), .Q(MVP1[7]), .QN(
        constructing_unit_Datapath_Last_register1_h_n51) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_h_MV_out_int_reg_8_ ( .D(
        constructing_unit_Datapath_Last_register1_h_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_h_n36), .Q(MVP1[8]), .QN(
        constructing_unit_Datapath_Last_register1_h_n50) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_h_MV_out_int_reg_9_ ( .D(
        constructing_unit_Datapath_Last_register1_h_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_h_n36), .Q(MVP1[9]), .QN(
        constructing_unit_Datapath_Last_register1_h_n49) );
  DFFR_X1 constructing_unit_Datapath_Last_register1_h_MV_out_int_reg_10_ ( .D(
        constructing_unit_Datapath_Last_register1_h_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register1_h_n36), .Q(MVP1[10]), .QN(
        constructing_unit_Datapath_Last_register1_h_n48) );
  INV_X1 constructing_unit_Datapath_Last_register2_h_U26 ( .A(
        constructing_unit_Datapath_n19), .ZN(
        constructing_unit_Datapath_Last_register2_h_n36) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_h_U25 ( .A1(
        constructing_unit_Datapath_MV2_int_h_13__9_), .A2(
        constructing_unit_Datapath_Last_register2_h_n33), .ZN(
        constructing_unit_Datapath_Last_register2_h_n60) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_h_U24 ( .B1(
        constructing_unit_Datapath_Last_register2_h_n49), .B2(
        constructing_unit_Datapath_Last_register2_h_n35), .A(
        constructing_unit_Datapath_Last_register2_h_n60), .ZN(
        constructing_unit_Datapath_Last_register2_h_n38) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_h_U23 ( .A1(
        constructing_unit_Datapath_MV2_int_h_13__8_), .A2(
        constructing_unit_Datapath_Last_register2_h_n33), .ZN(
        constructing_unit_Datapath_Last_register2_h_n61) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_h_U22 ( .B1(
        constructing_unit_Datapath_Last_register2_h_n50), .B2(
        constructing_unit_Datapath_Last_register2_h_n35), .A(
        constructing_unit_Datapath_Last_register2_h_n61), .ZN(
        constructing_unit_Datapath_Last_register2_h_n39) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_h_U21 ( .A1(
        constructing_unit_Datapath_MV2_int_h_13__7_), .A2(
        constructing_unit_Datapath_Last_register2_h_n33), .ZN(
        constructing_unit_Datapath_Last_register2_h_n62) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_h_U20 ( .B1(
        constructing_unit_Datapath_Last_register2_h_n51), .B2(
        constructing_unit_Datapath_Last_register2_h_n35), .A(
        constructing_unit_Datapath_Last_register2_h_n62), .ZN(
        constructing_unit_Datapath_Last_register2_h_n40) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_h_U19 ( .A1(
        constructing_unit_Datapath_MV2_int_h_13__6_), .A2(
        constructing_unit_Datapath_Last_register2_h_n33), .ZN(
        constructing_unit_Datapath_Last_register2_h_n63) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_h_U18 ( .B1(
        constructing_unit_Datapath_Last_register2_h_n52), .B2(
        constructing_unit_Datapath_Last_register2_h_n35), .A(
        constructing_unit_Datapath_Last_register2_h_n63), .ZN(
        constructing_unit_Datapath_Last_register2_h_n41) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_h_U17 ( .A1(
        constructing_unit_Datapath_MV2_int_h_13__5_), .A2(
        constructing_unit_Datapath_Last_register2_h_n33), .ZN(
        constructing_unit_Datapath_Last_register2_h_n64) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_h_U16 ( .B1(
        constructing_unit_Datapath_Last_register2_h_n53), .B2(
        constructing_unit_Datapath_Last_register2_h_n35), .A(
        constructing_unit_Datapath_Last_register2_h_n64), .ZN(
        constructing_unit_Datapath_Last_register2_h_n42) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_h_U15 ( .A1(
        constructing_unit_Datapath_MV2_int_h_13__4_), .A2(
        constructing_unit_Datapath_Last_register2_h_n33), .ZN(
        constructing_unit_Datapath_Last_register2_h_n65) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_h_U14 ( .B1(
        constructing_unit_Datapath_Last_register2_h_n54), .B2(
        constructing_unit_Datapath_Last_register2_h_n35), .A(
        constructing_unit_Datapath_Last_register2_h_n65), .ZN(
        constructing_unit_Datapath_Last_register2_h_n43) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_h_U13 ( .A1(
        constructing_unit_Datapath_MV2_int_h_13__3_), .A2(
        constructing_unit_Datapath_Last_register2_h_n33), .ZN(
        constructing_unit_Datapath_Last_register2_h_n66) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_h_U12 ( .B1(
        constructing_unit_Datapath_Last_register2_h_n55), .B2(
        constructing_unit_Datapath_Last_register2_h_n35), .A(
        constructing_unit_Datapath_Last_register2_h_n66), .ZN(
        constructing_unit_Datapath_Last_register2_h_n44) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_h_U11 ( .A1(
        constructing_unit_Datapath_MV2_int_h_13__2_), .A2(
        constructing_unit_Datapath_Last_register2_h_n33), .ZN(
        constructing_unit_Datapath_Last_register2_h_n67) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_h_U10 ( .B1(
        constructing_unit_Datapath_Last_register2_h_n56), .B2(
        constructing_unit_Datapath_Last_register2_h_n35), .A(
        constructing_unit_Datapath_Last_register2_h_n67), .ZN(
        constructing_unit_Datapath_Last_register2_h_n45) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_h_U9 ( .A1(
        constructing_unit_Datapath_MV2_int_h_13__1_), .A2(
        constructing_unit_Datapath_Last_register2_h_n33), .ZN(
        constructing_unit_Datapath_Last_register2_h_n68) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_h_U8 ( .B1(
        constructing_unit_Datapath_Last_register2_h_n57), .B2(
        constructing_unit_Datapath_Last_register2_h_n35), .A(
        constructing_unit_Datapath_Last_register2_h_n68), .ZN(
        constructing_unit_Datapath_Last_register2_h_n46) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_h_U7 ( .A1(
        constructing_unit_Datapath_MV2_int_h_13__0_), .A2(
        constructing_unit_Datapath_Last_register2_h_n33), .ZN(
        constructing_unit_Datapath_Last_register2_h_n69) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_h_U6 ( .B1(
        constructing_unit_Datapath_Last_register2_h_n58), .B2(
        constructing_unit_Datapath_Last_register2_h_n35), .A(
        constructing_unit_Datapath_Last_register2_h_n69), .ZN(
        constructing_unit_Datapath_Last_register2_h_n47) );
  NAND2_X1 constructing_unit_Datapath_Last_register2_h_U5 ( .A1(
        constructing_unit_Datapath_MV2_int_h_13__10_), .A2(
        constructing_unit_Datapath_Last_register2_h_n33), .ZN(
        constructing_unit_Datapath_Last_register2_h_n59) );
  OAI21_X1 constructing_unit_Datapath_Last_register2_h_U4 ( .B1(
        constructing_unit_Datapath_Last_register2_h_n48), .B2(
        constructing_unit_Datapath_Last_register2_h_n33), .A(
        constructing_unit_Datapath_Last_register2_h_n59), .ZN(
        constructing_unit_Datapath_Last_register2_h_n37) );
  BUF_X1 constructing_unit_Datapath_Last_register2_h_U3 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_Last_register2_h_n35) );
  BUF_X1 constructing_unit_Datapath_Last_register2_h_U2 ( .A(
        constructing_unit_Datapath_n1), .Z(
        constructing_unit_Datapath_Last_register2_h_n33) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_h_MV_out_int_reg_0_ ( .D(
        constructing_unit_Datapath_Last_register2_h_n47), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_h_n36), .Q(MVP2[0]), .QN(
        constructing_unit_Datapath_Last_register2_h_n58) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_h_MV_out_int_reg_1_ ( .D(
        constructing_unit_Datapath_Last_register2_h_n46), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_h_n36), .Q(MVP2[1]), .QN(
        constructing_unit_Datapath_Last_register2_h_n57) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_h_MV_out_int_reg_2_ ( .D(
        constructing_unit_Datapath_Last_register2_h_n45), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_h_n36), .Q(MVP2[2]), .QN(
        constructing_unit_Datapath_Last_register2_h_n56) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_h_MV_out_int_reg_3_ ( .D(
        constructing_unit_Datapath_Last_register2_h_n44), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_h_n36), .Q(MVP2[3]), .QN(
        constructing_unit_Datapath_Last_register2_h_n55) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_h_MV_out_int_reg_4_ ( .D(
        constructing_unit_Datapath_Last_register2_h_n43), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_h_n36), .Q(MVP2[4]), .QN(
        constructing_unit_Datapath_Last_register2_h_n54) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_h_MV_out_int_reg_5_ ( .D(
        constructing_unit_Datapath_Last_register2_h_n42), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_h_n36), .Q(MVP2[5]), .QN(
        constructing_unit_Datapath_Last_register2_h_n53) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_h_MV_out_int_reg_6_ ( .D(
        constructing_unit_Datapath_Last_register2_h_n41), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_h_n36), .Q(MVP2[6]), .QN(
        constructing_unit_Datapath_Last_register2_h_n52) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_h_MV_out_int_reg_7_ ( .D(
        constructing_unit_Datapath_Last_register2_h_n40), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_h_n36), .Q(MVP2[7]), .QN(
        constructing_unit_Datapath_Last_register2_h_n51) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_h_MV_out_int_reg_8_ ( .D(
        constructing_unit_Datapath_Last_register2_h_n39), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_h_n36), .Q(MVP2[8]), .QN(
        constructing_unit_Datapath_Last_register2_h_n50) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_h_MV_out_int_reg_9_ ( .D(
        constructing_unit_Datapath_Last_register2_h_n38), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_h_n36), .Q(MVP2[9]), .QN(
        constructing_unit_Datapath_Last_register2_h_n49) );
  DFFR_X1 constructing_unit_Datapath_Last_register2_h_MV_out_int_reg_10_ ( .D(
        constructing_unit_Datapath_Last_register2_h_n37), .CK(clk), .RN(
        constructing_unit_Datapath_Last_register2_h_n36), .Q(MVP2[10]), .QN(
        constructing_unit_Datapath_Last_register2_h_n48) );
  OR2_X1 extimating_unit_U2 ( .A1(cDONE), .A2(VALID), .ZN(
        extimating_unit_VALID_int) );
  AND2_X1 extimating_unit_U1 ( .A1(eREADY), .A2(extimating_unit_VALID_int), 
        .ZN(extimating_unit_RF_in_WE_int) );
  CLKBUF_X3 extimating_unit_Pixel_Retrieval_Unit_U166 ( .A(
        extimating_unit_RST2_int), .Z(extimating_unit_Pixel_Retrieval_Unit_n36) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U164 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_block_num[1]), .A2(extimating_unit_Pixel_Retrieval_Unit_n21), .B1(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_block_num[1]), .B2(extimating_unit_Pixel_Retrieval_Unit_n19), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n97) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U163 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n97), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n129) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U162 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_CurCU_h_short_0_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n21), .B1(
        extimating_unit_Pixel_Retrieval_Unit_CurCU_w_short_0_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n19), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n98) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U161 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n98), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n130) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U160 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__11_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n39) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U159 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__5_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n51) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U158 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n53) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U157 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__3_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n55) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U156 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__10_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n41) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U155 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__9_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n43) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U154 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__8_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n45) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U153 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__7_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n47) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U152 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n49) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U151 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[9]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n42) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U150 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n43), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n30), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n42), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[33]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U149 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[8]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n44) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U148 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n45), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n30), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n44), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[32]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U147 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[7]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n46) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U146 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n47), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n30), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n46), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[31]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U145 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[6]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n48) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U144 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n49), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n29), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n48), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[30]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U143 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[5]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n50) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U142 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n51), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n29), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n50), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[29]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U141 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[4]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n52) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U140 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n53), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n31), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n52), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[28]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U139 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[3]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n54) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U138 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n55), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n30), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n54), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[27]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U137 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[2]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n56) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U136 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n57), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n32), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n56), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[26]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U135 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[1]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n58) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U134 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n59), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n31), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n58), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[25]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U133 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n60), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n31), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n60), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[24]) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U132 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sixPar_samp), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n17) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U131 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sixPar_samp), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n16) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_U130 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n5), .A2(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n9) );
  XNOR2_X1 extimating_unit_Pixel_Retrieval_Unit_U129 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__5_), .B(
        extimating_unit_Pixel_Retrieval_Unit_n9), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n8) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_U128 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__4_), .B(
        extimating_unit_Pixel_Retrieval_Unit_n5), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n7) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_U127 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__2_), .B(
        extimating_unit_Pixel_Retrieval_Unit_add_239_carry_2_), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U126 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__2_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n57) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U125 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n59) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_U124 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n4), .A2(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__3_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n5) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_U123 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_add_239_carry_2_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__2_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n4) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_U122 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_y_count_out_0_), .B(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__0_), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n3) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U121 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n60) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U120 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[10]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n40) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U119 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n41), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n31), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[34]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U118 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n38) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U117 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n39), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n32), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[35]) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_U116 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__0_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_y_count_out_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n2) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_U115 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__3_), .B(
        extimating_unit_Pixel_Retrieval_Unit_n4), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n1) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U114 ( .A1(
        extimating_unit_MV1_out_int[10]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_MV2_out_int[21]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n84) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U113 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n84), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n61) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U112 ( .A1(
        extimating_unit_MV1_out_int[21]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B1(
        extimating_unit_MV2_out_int[10]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n26), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n95) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U111 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n95), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n118) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U110 ( .A(
        extimating_unit_MV0_out_int[10]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n72) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U109 ( .A(
        extimating_unit_MV0_out_int[21]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n107) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U108 ( .A(
        extimating_unit_MV0_out_int[20]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n108) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U107 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n17), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n11) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U106 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n17), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n12) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U105 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n16), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n15) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U104 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n16), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n13) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U103 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n16), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n14) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U102 ( .A1(
        extimating_unit_MV1_out_int[11]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B1(
        extimating_unit_MV2_out_int[0]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n26), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n96) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U101 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n96), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n128) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U100 ( .A1(
        extimating_unit_MV1_out_int[0]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_MV2_out_int[11]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n85) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U99 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n85), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n71) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U98 ( .A1(
        extimating_unit_MV1_out_int[9]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n35), .B2(
        extimating_unit_MV2_out_int[20]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n75) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U97 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n62) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U96 ( .A1(
        extimating_unit_MV1_out_int[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_MV2_out_int[19]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n21), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n76) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U95 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n76), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n63) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U94 ( .A1(
        extimating_unit_MV1_out_int[7]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_MV2_out_int[18]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n22), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n77) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U93 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n77), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n64) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U92 ( .A1(
        extimating_unit_MV1_out_int[6]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_MV2_out_int[17]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n21), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n78) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U91 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n78), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n65) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U90 ( .A1(
        extimating_unit_MV1_out_int[5]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_MV2_out_int[16]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n22), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n79) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U89 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n79), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n66) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U88 ( .A1(
        extimating_unit_MV1_out_int[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_MV2_out_int[15]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n22), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n80) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U87 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n80), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n67) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U86 ( .A1(
        extimating_unit_MV1_out_int[3]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_MV2_out_int[14]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n22), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n81) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U85 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n81), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n68) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U84 ( .A1(
        extimating_unit_MV1_out_int[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_MV2_out_int[13]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n82) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U83 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n82), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n69) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U82 ( .A1(
        extimating_unit_MV1_out_int[20]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B1(
        extimating_unit_MV2_out_int[9]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n24), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n86) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U81 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n86), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n119) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U80 ( .A1(
        extimating_unit_MV1_out_int[19]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B1(
        extimating_unit_MV2_out_int[8]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n24), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n87) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U79 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n87), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n120) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U78 ( .A1(
        extimating_unit_MV1_out_int[18]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_MV2_out_int[7]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n24), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n88) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U77 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n88), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n121) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U76 ( .A1(
        extimating_unit_MV1_out_int[17]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B1(
        extimating_unit_MV2_out_int[6]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n24), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n89) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U75 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n89), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n122) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U74 ( .A1(
        extimating_unit_MV1_out_int[16]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B1(
        extimating_unit_MV2_out_int[5]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n25), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n90) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U73 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n90), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n123) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U72 ( .A1(
        extimating_unit_MV1_out_int[15]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B1(
        extimating_unit_MV2_out_int[4]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n25), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n91) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U71 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n91), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n124) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U70 ( .A1(
        extimating_unit_MV1_out_int[14]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B1(
        extimating_unit_MV2_out_int[3]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n25), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n92) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U69 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n92), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n125) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U68 ( .A1(
        extimating_unit_MV1_out_int[13]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B1(
        extimating_unit_MV2_out_int[2]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n25), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n93) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U67 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n93), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n126) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U66 ( .A(
        extimating_unit_MV0_out_int[9]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n73) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U65 ( .A(
        extimating_unit_MV0_out_int[8]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n74) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U64 ( .A(
        extimating_unit_MV0_out_int[7]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n99) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U63 ( .A(
        extimating_unit_MV0_out_int[6]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n100) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U62 ( .A(
        extimating_unit_MV0_out_int[5]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n101) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U61 ( .A(
        extimating_unit_MV0_out_int[4]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n102) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U60 ( .A(
        extimating_unit_MV0_out_int[3]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n103) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U59 ( .A(
        extimating_unit_MV0_out_int[2]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n104) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U58 ( .A(
        extimating_unit_MV0_out_int[1]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n105) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U57 ( .A(
        extimating_unit_MV0_out_int[19]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n109) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U56 ( .A(
        extimating_unit_MV0_out_int[18]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n110) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U55 ( .A(
        extimating_unit_MV0_out_int[17]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n111) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U54 ( .A(
        extimating_unit_MV0_out_int[16]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n112) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U53 ( .A(
        extimating_unit_MV0_out_int[15]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n113) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U52 ( .A(
        extimating_unit_MV0_out_int[14]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n114) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U51 ( .A(
        extimating_unit_MV0_out_int[13]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n115) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U50 ( .A(
        extimating_unit_MV0_out_int[12]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n116) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U49 ( .A(
        extimating_unit_MV0_out_int[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n106) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U48 ( .A(
        extimating_unit_MV0_out_int[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n117) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U47 ( .A1(
        extimating_unit_MV1_out_int[12]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B1(
        extimating_unit_MV2_out_int[1]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n26), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n94) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_U46 ( .A1(
        extimating_unit_MV1_out_int[1]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B1(
        extimating_unit_MV2_out_int[12]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n83) );
  BUF_X2 extimating_unit_Pixel_Retrieval_Unit_U45 ( .A(
        extimating_unit_RST2_int), .Z(extimating_unit_Pixel_Retrieval_Unit_n37) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U44 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n34), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n107), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n72), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__10_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U43 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n19), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n107), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n29), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n72), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__10_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U42 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n83), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n70) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U41 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n15), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n35) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U40 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n33), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n117), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n106), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__0_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U39 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n117), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n29), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n106), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__0_) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U38 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n15), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n34) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U37 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n15), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n33) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U36 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n14), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n32) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U35 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n94), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n127) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U34 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n12), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n26) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U33 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n11), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n22) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U32 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n11), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n23) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U31 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n12), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n24) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U30 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n12), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n25) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U29 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n11), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n21) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U28 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n13), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n28) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U27 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n14), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n31) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n14), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n30) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U25 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n13), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n29) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_U24 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n13), .Z(
        extimating_unit_Pixel_Retrieval_Unit_n27) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U23 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n108), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n26), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n73), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__9_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U22 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n109), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n27), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n74), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__8_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U21 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n110), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n27), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n99), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__7_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U20 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n111), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n27), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n100), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__6_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U19 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n112), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n27), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n101), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__5_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U18 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n113), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n28), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n102), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__4_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U17 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n114), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n28), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n103), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__3_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U16 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n115), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n28), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n104), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__2_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U15 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n116), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n28), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n105), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__1_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U14 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n32), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n108), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n73), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__9_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U13 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n34), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n109), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n18), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n74), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__8_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U12 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n34), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n110), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n19), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n99), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__7_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U11 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n33), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n111), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n100), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__6_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U10 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n32), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n112), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n101), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__5_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U9 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n34), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n113), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n102), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__4_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U8 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n33), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n114), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n103), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__3_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U7 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n35), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n115), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n104), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__2_) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_U6 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n33), .A2(
        extimating_unit_Pixel_Retrieval_Unit_n116), .B1(
        extimating_unit_Pixel_Retrieval_Unit_n20), .B2(
        extimating_unit_Pixel_Retrieval_Unit_n105), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__1_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n31), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n20) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n28), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n19) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n27), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_n18) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_add_239_U1_1 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__1_), .B(
        extimating_unit_Pixel_Retrieval_Unit_y_count_out_1_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_n2), .CO(
        extimating_unit_Pixel_Retrieval_Unit_add_239_carry_2_), .S(
        extimating_unit_Pixel_Retrieval_Unit_y_short_1_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_width_register_U3 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_width_register_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_width_register_Q_int_reg_0_ ( 
        .D(CU_w[5]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_width_register_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_CurCU_w_short_0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_width_register_Q_int_reg_1_ ( 
        .D(CU_w[6]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_width_register_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_block_num[1]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_height_register_U3 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_height_register_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_height_register_Q_int_reg_0_ ( 
        .D(CU_h[5]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_height_register_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_CurCU_h_short_0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_height_register_Q_int_reg_1_ ( 
        .D(CU_h[6]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_height_register_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_block_num[1]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_sixPar_reg_U3 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sixPar_reg_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_sixPar_reg_Q_int_reg ( .D(
        sixPar), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_sixPar_reg_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sixPar_samp) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U351 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n94), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n83), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n69), .ZN(
        extimating_unit_MV2_out_int[10]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U350 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n93), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n82), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n69), .ZN(
        extimating_unit_MV2_out_int[9]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U349 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n92), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n81), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n69), .ZN(
        extimating_unit_MV2_out_int[8]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U348 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n204), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n193), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n347), .ZN(
        extimating_unit_MV2_out_int[21]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U347 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n203), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n192), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n347), .ZN(
        extimating_unit_MV2_out_int[20]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U346 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n115), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n104), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n72), .ZN(
        extimating_unit_MV1_out_int[20]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U345 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n137), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n126), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n338), .ZN(
        extimating_unit_MV1_out_int[9]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U344 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n160), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n149), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n341), .ZN(
        extimating_unit_MV0_out_int[21]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U343 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n159), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n148), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n341), .ZN(
        extimating_unit_MV0_out_int[20]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U342 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n182), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n171), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n344), .ZN(
        extimating_unit_MV0_out_int[10]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U341 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n116), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n105), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n72), .ZN(
        extimating_unit_MV1_out_int[21]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U340 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n138), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n127), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n339), .ZN(
        extimating_unit_MV1_out_int[10]) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U339 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_samp), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n63) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U338 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_samp), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n62) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U337 ( .A(n233), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n404) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U336 ( .A(n234), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n405) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U335 ( .A(n235), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n406) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U334 ( .A(n236), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n407) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U333 ( .A(n237), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n408) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U332 ( .A(n238), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n409) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U331 ( .A(n239), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n410) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U330 ( .A(n240), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n411) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U329 ( .A(n241), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n412) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U328 ( .A(n242), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n413) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U327 ( .A(n243), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n414) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U326 ( .A(n201), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n372) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U325 ( .A(n202), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n373) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U324 ( .A(n203), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n374) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U323 ( .A(n204), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n375) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U322 ( .A(n205), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n376) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U321 ( .A(n206), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n377) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U320 ( .A(n200), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n371) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U319 ( .A(n207), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n378) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U318 ( .A(n208), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n379) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U317 ( .A(n209), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n380) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U316 ( .A(n210), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n381) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U315 ( .A(n190), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n361) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U314 ( .A(n191), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n362) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U313 ( .A(n192), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n363) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U312 ( .A(n193), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n364) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U311 ( .A(n194), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n365) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U310 ( .A(n195), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n366) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U309 ( .A(n196), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n367) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U308 ( .A(n197), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n368) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U307 ( .A(n211), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n382) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U306 ( .A(n212), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n383) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U305 ( .A(n213), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n384) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U304 ( .A(n214), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n385) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U303 ( .A(n215), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n386) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U302 ( .A(n216), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n387) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U301 ( .A(n217), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n388) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U300 ( .A(n218), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n389) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U299 ( .A(n219), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n390) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U298 ( .A(n220), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n391) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U297 ( .A(n221), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n392) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U296 ( .A(n178), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n349) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U295 ( .A(n179), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n350) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U294 ( .A(n180), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n351) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U293 ( .A(n181), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n352) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U292 ( .A(n182), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n353) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U291 ( .A(n183), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n354) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U290 ( .A(n184), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n355) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U289 ( .A(n185), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n356) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U288 ( .A(n186), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n357) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U287 ( .A(n187), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n358) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U286 ( .A(n188), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n359) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U285 ( .A(n222), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n393) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U284 ( .A(n223), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n394) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U283 ( .A(n224), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n395) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U282 ( .A(n225), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n396) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U281 ( .A(n226), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n397) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U280 ( .A(n227), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n398) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U279 ( .A(n228), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n399) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U278 ( .A(n229), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n400) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U277 ( .A(n230), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n401) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U276 ( .A(n231), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n402) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U275 ( .A(n232), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n403) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U274 ( .A(n189), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n360) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U273 ( .A(n198), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n369) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U272 ( .A(n199), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n370) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U271 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n17), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n377), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n198), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n330) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U270 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n18), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n378), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n197), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n329) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U269 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n18), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n379), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n196), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n328) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U268 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n18), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n380), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n195), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n327) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U267 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n19), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n381), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n194), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n326) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U266 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n19), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n382), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n182), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n314) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U265 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n19), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n383), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n181), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n313) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U264 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n19), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n384), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n180), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n312) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U263 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n385), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n179), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n311) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U262 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n386), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n178), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n310) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U261 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n387), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n177), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n309) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U260 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n20), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n388), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n176), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n308) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U259 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n24), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n371), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n204), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n337) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U258 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n18), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n372), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n203), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n335) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U257 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n17), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n373), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n202), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n334) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U256 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n16), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n374), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n201), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n333) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U255 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n17), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n375), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n200), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n332) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U254 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n17), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n376), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n199), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n331) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U253 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n42), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n371), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n193), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n325) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U252 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n42), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n372), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n192), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n324) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U251 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n42), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n373), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n191), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n323) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U250 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n42), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n374), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n190), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n322) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U249 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n42), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n375), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n189), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n321) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U248 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n43), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n376), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n188), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n320) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U247 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n21), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n389), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n175), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n307) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U246 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n21), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n390), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n174), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n306) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U245 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n21), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n391), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n173), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n305) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U244 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n21), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n392), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n172), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n304) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U243 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n22), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n349), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n160), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n292) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U242 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n22), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n350), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n159), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n291) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U241 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n22), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n351), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n158), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n290) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U240 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n22), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n352), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n157), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n289) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U239 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n23), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n353), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n156), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n288) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U238 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n23), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n354), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n155), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n287) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U237 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n23), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n355), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n154), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n286) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U236 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n23), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n356), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n153), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n285) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U235 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n24), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n357), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n152), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n284) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U234 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n24), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n358), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n151), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n283) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U233 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n24), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n359), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n150), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n282) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U232 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n25), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n393), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n138), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n270) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U231 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n25), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n394), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n137), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n269) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U230 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n25), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n395), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n136), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n268) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U229 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n25), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n396), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n135), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n267) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U228 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n26), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n397), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n134), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n266) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U227 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n26), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n398), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n133), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n265) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U226 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n26), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n399), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n132), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n264) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U225 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n26), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n400), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n131), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n263) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U224 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n27), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n401), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n130), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n262) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U223 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n27), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n402), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n129), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n261) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U222 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n27), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n403), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n128), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n260) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U221 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n27), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n360), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n116), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n248) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U220 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n28), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n361), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n115), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n247) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U219 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n28), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n362), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n114), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n246) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U218 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n28), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n363), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n113), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n245) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U217 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n28), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n364), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n112), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n244) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U216 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n29), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n365), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n111), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n243) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U215 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n29), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n366), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n110), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n242) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U214 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n29), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n367), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n109), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n241) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U213 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n29), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n368), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n108), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n240) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U212 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n30), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n369), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n107), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n239) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U211 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n30), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n370), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n106), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n238) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U210 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n404), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n15), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n94), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n226) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U209 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n405), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n16), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n93), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n225) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U208 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n406), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n16), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n92), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n224) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U207 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n407), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n15), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n91), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n223) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U206 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n408), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n16), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n90), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n222) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U205 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n409), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n15), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n89), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n221) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U204 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n410), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n13), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n88), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n220) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U203 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n411), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n15), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n87), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n219) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U202 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n412), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n13), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n86), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n218) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U201 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n413), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n13), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n85), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n217) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U200 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n414), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n13), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n84), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n216) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U199 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n43), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n377), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n187), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n319) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U198 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n43), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n378), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n186), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n318) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U197 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n43), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n379), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n185), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n317) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U196 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n43), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n380), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n184), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n316) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U195 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n44), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n381), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n183), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n315) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U194 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n44), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n382), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n171), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n303) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U193 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n44), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n383), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n170), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n302) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U192 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n44), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n384), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n169), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n301) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U191 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n44), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n385), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n168), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n300) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U190 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n45), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n386), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n167), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n299) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U189 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n45), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n387), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n166), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n298) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U188 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n45), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n388), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n165), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n297) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U187 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n45), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n389), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n164), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n296) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U186 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n45), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n390), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n163), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n295) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U185 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n46), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n391), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n162), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n294) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U184 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n46), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n392), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n161), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n293) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U183 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n46), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n349), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n149), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n281) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U182 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n46), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n350), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n148), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n280) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U181 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n46), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n351), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n147), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n279) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U180 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n47), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n352), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n146), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n278) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U179 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n47), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n353), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n145), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n277) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U178 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n47), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n354), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n144), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n276) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U177 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n47), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n355), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n143), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n275) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U176 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n47), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n356), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n274) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U175 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n48), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n357), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n141), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n273) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U174 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n48), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n358), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n140), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n272) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U173 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n48), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n359), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n139), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n271) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U172 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n48), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n393), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n127), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n259) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U171 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n48), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n394), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n126), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n258) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U170 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n49), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n395), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n125), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n257) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U169 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n49), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n396), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n124), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n256) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U168 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n49), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n397), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n123), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n255) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U167 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n49), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n398), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n122), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n254) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U166 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n49), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n399), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n121), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n253) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U165 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n50), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n400), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n120), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n252) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U164 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n50), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n401), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n119), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n251) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U163 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n50), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n402), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n118), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n250) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U162 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n50), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n403), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n117), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n249) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U161 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n50), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n360), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n105), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n237) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U160 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n51), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n361), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n104), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n236) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U159 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n51), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n362), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n103), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n235) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U158 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n51), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n363), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n102), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n234) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U157 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n51), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n364), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n101), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n233) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U156 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n51), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n365), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n100), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n232) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U155 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n52), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n366), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n99), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n231) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U154 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n52), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n367), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n98), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n230) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U153 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n52), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n368), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n97), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n229) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U152 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n52), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n369), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n96), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n228) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U151 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n52), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n370), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n95), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n227) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U150 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n53), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n404), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n83), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n215) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U149 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n53), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n405), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n82), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n214) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U148 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n53), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n406), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n81), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n213) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U147 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n53), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n407), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n80), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n212) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U146 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n53), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n408), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n79), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n211) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U145 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n54), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n409), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n78), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n210) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U144 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n54), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n410), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n77), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n209) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U143 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n54), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n411), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n76), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n208) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U142 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n54), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n412), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n75), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n207) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U141 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n54), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n413), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n74), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n206) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U140 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n55), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n414), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n73), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n205) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U139 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n202), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n191), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n346), .ZN(
        extimating_unit_MV2_out_int[19]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U138 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n201), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n190), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n346), .ZN(
        extimating_unit_MV2_out_int[18]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U137 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n200), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n189), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n346), .ZN(
        extimating_unit_MV2_out_int[17]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U136 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n199), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n188), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n346), .ZN(
        extimating_unit_MV2_out_int[16]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U135 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n198), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n187), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n345), .ZN(
        extimating_unit_MV2_out_int[15]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U134 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n197), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n186), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n345), .ZN(
        extimating_unit_MV2_out_int[14]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U133 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n196), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n185), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n345), .ZN(
        extimating_unit_MV2_out_int[13]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U132 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n195), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n184), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n345), .ZN(
        extimating_unit_MV2_out_int[12]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U131 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n91), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n80), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n68), .ZN(
        extimating_unit_MV2_out_int[7]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U130 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n90), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n79), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n68), .ZN(
        extimating_unit_MV2_out_int[6]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U129 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n89), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n78), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n68), .ZN(
        extimating_unit_MV2_out_int[5]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U128 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n88), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n77), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n68), .ZN(
        extimating_unit_MV2_out_int[4]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U127 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n87), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n76), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n67), .ZN(
        extimating_unit_MV2_out_int[3]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U126 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n86), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n75), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n67), .ZN(
        extimating_unit_MV2_out_int[2]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U125 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n85), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n74), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n67), .ZN(
        extimating_unit_MV2_out_int[1]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U124 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n194), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n183), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n344), .ZN(
        extimating_unit_MV2_out_int[11]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U123 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n84), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n73), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n67), .ZN(
        extimating_unit_MV2_out_int[0]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U122 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n114), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n103), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n71), .ZN(
        extimating_unit_MV1_out_int[19]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U121 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n113), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n102), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n71), .ZN(
        extimating_unit_MV1_out_int[18]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U120 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n112), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n101), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n71), .ZN(
        extimating_unit_MV1_out_int[17]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U119 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n111), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n100), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n71), .ZN(
        extimating_unit_MV1_out_int[16]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U118 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n110), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n99), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n70), .ZN(
        extimating_unit_MV1_out_int[15]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U117 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n109), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n98), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n70), .ZN(
        extimating_unit_MV1_out_int[14]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U116 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n108), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n97), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n70), .ZN(
        extimating_unit_MV1_out_int[13]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U115 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n107), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n96), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n70), .ZN(
        extimating_unit_MV1_out_int[12]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U114 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n136), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n125), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n338), .ZN(
        extimating_unit_MV1_out_int[8]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U113 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n135), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n124), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n338), .ZN(
        extimating_unit_MV1_out_int[7]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U112 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n134), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n123), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n338), .ZN(
        extimating_unit_MV1_out_int[6]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U111 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n133), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n122), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n336), .ZN(
        extimating_unit_MV1_out_int[5]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U110 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n132), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n121), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n336), .ZN(
        extimating_unit_MV1_out_int[4]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U109 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n131), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n120), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n336), .ZN(
        extimating_unit_MV1_out_int[3]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U108 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n130), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n119), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n336), .ZN(
        extimating_unit_MV1_out_int[2]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U107 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n129), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n118), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n72), .ZN(
        extimating_unit_MV1_out_int[1]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U106 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n158), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n147), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n341), .ZN(
        extimating_unit_MV0_out_int[19]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U105 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n157), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n146), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n341), .ZN(
        extimating_unit_MV0_out_int[18]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U104 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n156), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n145), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n340), .ZN(
        extimating_unit_MV0_out_int[17]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U103 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n155), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n144), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n340), .ZN(
        extimating_unit_MV0_out_int[16]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U102 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n154), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n143), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n340), .ZN(
        extimating_unit_MV0_out_int[15]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U101 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n153), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n340), .ZN(
        extimating_unit_MV0_out_int[14]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U100 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n152), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n141), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n339), .ZN(
        extimating_unit_MV0_out_int[13]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U99 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n151), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n140), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n339), .ZN(
        extimating_unit_MV0_out_int[12]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U98 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n181), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n170), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n344), .ZN(
        extimating_unit_MV0_out_int[9]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U97 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n180), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n169), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n344), .ZN(
        extimating_unit_MV0_out_int[8]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U96 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n168), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n343), .ZN(
        extimating_unit_MV0_out_int[7]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U95 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n178), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n167), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n343), .ZN(
        extimating_unit_MV0_out_int[6]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U94 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n177), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n166), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n343), .ZN(
        extimating_unit_MV0_out_int[5]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U93 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n165), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n343), .ZN(
        extimating_unit_MV0_out_int[4]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U92 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n175), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n164), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n342), .ZN(
        extimating_unit_MV0_out_int[3]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U91 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n174), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n163), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n342), .ZN(
        extimating_unit_MV0_out_int[2]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U90 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n162), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n342), .ZN(
        extimating_unit_MV0_out_int[1]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U89 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n150), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n139), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n339), .ZN(
        extimating_unit_MV0_out_int[11]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U88 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n172), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n161), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n342), .ZN(
        extimating_unit_MV0_out_int[0]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U87 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n106), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n95), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n69), .ZN(
        extimating_unit_MV1_out_int[11]) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U86 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n128), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65), .B1(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n117), .B2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n72), .ZN(
        extimating_unit_MV1_out_int[0]) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U85 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n63), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n57) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U84 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n62), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n59) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U83 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n63), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n58) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U82 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n63), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n56) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U81 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n62), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n60) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U80 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n62), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n61) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U79 ( .A(
        extimating_unit_RF_Addr_DP_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n415) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U78 ( .A1(
        extimating_unit_RF_in_WE_int), .A2(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n415), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n1) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U77 ( .A1(
        extimating_unit_RF_Addr_DP_int), .A2(extimating_unit_RF_in_WE_int), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_input_RF_n14) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U76 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n38) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U75 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n14), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n8) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U74 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n14), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n9) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U73 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n37) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U72 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n61), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n348) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U71 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n57), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n72) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U70 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n57), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n71) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U69 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n57), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n70) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U68 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n58), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n338) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U67 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n58), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n336) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U66 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n59), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n341) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U65 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n59), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n340) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U64 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n58), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n339) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U63 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n60), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n343) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U62 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n59), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n342) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U61 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n61), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n346) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U60 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n60), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n345) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U59 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n56), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n69) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U58 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n56), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n68) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U57 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n56), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n67) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U56 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n60), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n344) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U55 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n61), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n347) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U54 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n37), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n36) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U53 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n38), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n32) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U52 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n38), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n33) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U51 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n8), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n5) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U50 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n9), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n3) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U49 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n9), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n2) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U48 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n9), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n4) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U47 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n37), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n34) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U46 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n8), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n6) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U45 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n37), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n35) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U44 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n8), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U43 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n348), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n66) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U42 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n347), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n65) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U41 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n347), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n64) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U40 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n7), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n31) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U39 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n5), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n24) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U38 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n3), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n18) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U37 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n3), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n17) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U36 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n3), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n19) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U35 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n4), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n20) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U34 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n4), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n21) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U33 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n4), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n22) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U32 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n5), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n23) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U31 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n5), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n25) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U30 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n6), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n26) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U29 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n6), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n27) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U28 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n6), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n28) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U27 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n7), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n29) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n2), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n16) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U25 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n2), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n15) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U24 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n2), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n13) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U23 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n36), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n54) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U22 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n32), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n42) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U21 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n32), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n43) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U20 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n32), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n44) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U19 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n33), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n45) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U18 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n33), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n46) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U17 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n33), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n47) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U16 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n34), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n48) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U15 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n34), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n49) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U14 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n34), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n50) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n35), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n51) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U12 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n35), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n52) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n35), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n53) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n7), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n30) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n36), .Z(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n55) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n31), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n12) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n30), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n11) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U6 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n30), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n10) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n41) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n40) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n39) );
  INV_X8 extimating_unit_Pixel_Retrieval_Unit_input_RF_U2 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_0__0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n293), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n161) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_0__1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n294), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n162) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_0__2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n295), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n163) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_0__3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n296), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n164) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_0__4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n297), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n165) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_0__5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n298), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n166) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_0__6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n299), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n167) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_0__7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n300), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n168) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_0__8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n301), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n169) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_0__9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n302), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n170) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_0__10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n303), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n171) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_0__0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n271), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n139) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_0__1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n272), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n140) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_0__2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n273), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n141) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_0__3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n274), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n142) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_0__4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n275), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n143) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_0__5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n276), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n144) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_0__6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n277), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n145) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_0__7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n278), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n146) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_0__8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n279), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n147) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_0__9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n280), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n148) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_0__10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n281), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n149) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_0__0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n249), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n117) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_0__1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n250), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n118) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_0__2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n251), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n119) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_0__3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n252), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n120) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_0__4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n253), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n121) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_0__5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n254), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n122) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_0__6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n255), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n123) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_0__7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n256), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n124) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_0__8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n257), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n125) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_0__9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n258), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n126) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_0__10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n259), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n127) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_0__0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n227), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n95) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_0__1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n228), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n96) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_0__2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n229), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n97) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_0__3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n230), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n98) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_0__4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n231), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n99) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_0__5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n232), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n100) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_0__6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n233), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n101) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_0__7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n234), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n102) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_0__8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n235), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n103) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_0__9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n236), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n104) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_0__10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n237), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n105) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_0__0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n205), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n73) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_0__1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n206), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n74) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_0__2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n207), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n75) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_0__3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n208), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n76) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_0__4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n209), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n77) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_0__5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n210), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n78) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_0__6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n211), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n79) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_0__7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n212), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n80) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_0__8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n213), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n81) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_0__9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n214), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n82) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_0__10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n215), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n83) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_0__0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n315), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n183) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_0__1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n316), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n184) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_0__2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n317), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n185) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_0__3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n318), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n186) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_0__4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n319), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n187) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_1__0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n304), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n172) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_1__1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n305), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n173) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_1__2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n306), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n174) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_1__3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n307), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n175) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_1__0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n282), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n150) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_1__1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n283), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n151) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_1__2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n284), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n152) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_1__3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n285), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n153) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_1__4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n286), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n154) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_1__5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n287), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n155) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_1__6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n288), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n156) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_1__7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n289), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n157) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_1__8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n290), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n158) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_1__9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n291), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n159) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_v_reg_1__10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n292), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n160) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_1__0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n260), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n128) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_1__1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n261), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n129) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_1__2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n262), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n130) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_1__3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n263), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n131) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_1__4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n264), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n132) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_1__5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n265), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n133) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_1__6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n266), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n134) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_1__7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n267), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n135) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_1__8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n268), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n136) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_1__9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n269), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n137) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_h_reg_1__10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n270), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n138) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_1__0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n238), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n106) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_1__1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n239), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n107) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_1__2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n240), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n108) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_1__3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n241), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n109) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_1__4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n242), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n110) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_1__5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n243), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n111) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_1__6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n244), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n112) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_1__7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n245), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n113) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_1__8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n246), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n114) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_1__9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n247), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n115) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV1_v_reg_1__10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n248), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n116) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_1__0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n216), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n84) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_1__1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n217), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n85) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_1__2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n218), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n86) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_1__3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n219), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n87) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_1__4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n220), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n88) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_1__5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n221), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n89) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_1__6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n222), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n90) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_1__7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n223), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n91) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_1__8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n224), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n92) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_1__9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n225), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n93) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_h_reg_1__10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n226), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n94) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_0__5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n320), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n188) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_0__6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n321), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n189) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_0__7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n322), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n190) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_0__8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n323), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n191) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_0__9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n324), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n192) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_0__10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n325), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n193) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_1__4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n308), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n176) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_1__5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n309), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n177) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_1__6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n310), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n178) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_1__7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n311), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n179) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_1__8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n312), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n180) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_1__9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n313), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n181) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV0_h_reg_1__10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n314), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n182) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_1__0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n326), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n194) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_1__1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n327), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n195) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_1__2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n328), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n196) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_1__3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n329), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n197) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_1__4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n330), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n198) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_1__5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n331), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n199) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_1__6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n332), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n200) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_1__7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n333), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n201) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_1__8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n334), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n202) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_1__9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n335), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n203) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_MV2_v_reg_1__10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n337), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n416), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_n204) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_U4 ( 
        .A1(1'b1), .A2(extimating_unit_RF_Addr_DP_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_n7) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_U3 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_n6), 
        .B2(1'b1), .A(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_n7), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_n5)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_U2 ( 
        .A(extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_n3) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_n5), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_n3), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_samp), .QN(
        extimating_unit_Pixel_Retrieval_Unit_input_RF_RF_Addr_sampling_n6) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_U3 ( 
        .A1(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_n1), .A2(extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_n2), 
        .ZN(last_block_x) );
  OR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_U2 ( 
        .A1(extimating_unit_RST1_int), .A2(extimating_unit_RST_BLKx_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_count_RST) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_U5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_x0_int_0__5_), .B(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_block_num[1]), .Z(extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_n1)
         );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_U4 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_x0_int_0__4_), .B(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_block_num[0]), .Z(extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_n2)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurRep_U2 ( 
        .A(extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurRep_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurRep_tmp_reg ( 
        .D(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurRep_n2), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurRep_n1), .Q(extimating_unit_Pixel_Retrieval_Unit_x0_int_0__3_) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurRep_U3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_x0_int_0__3_), .B(
        extimating_unit_CE_REPx_int), .Z(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurRep_n2) );
  XNOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_U6 ( 
        .A(extimating_unit_CE_BLKx_int), .B(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_0__4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n3) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_U5 ( 
        .A1(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_count_RST), .A2(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n3), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n5) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_U4 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_x0_int_0__4_), .A2(
        extimating_unit_CE_BLKx_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n2) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_U3 ( 
        .A1(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_count_RST), .A2(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n4) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_U7 ( 
        .A(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n2), .B(extimating_unit_Pixel_Retrieval_Unit_x0_int_0__5_), .Z(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n1) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_count_tmp_reg_1_ ( 
        .D(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n4), .CK(clk), .Q(extimating_unit_Pixel_Retrieval_Unit_x0_int_0__5_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_count_tmp_reg_0_ ( 
        .D(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_CurBlock_n5), .CK(clk), .Q(extimating_unit_Pixel_Retrieval_Unit_x0_int_0__4_) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_encoder_U1 ( 
        .A(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_block_num[1]), .B(extimating_unit_Pixel_Retrieval_Unit_CurCU_w_short_0_), .Z(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_block_num[0]) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_U3 ( 
        .A1(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_n4), .A2(extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_n3), 
        .ZN(last_block_y) );
  OR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_U2 ( 
        .A1(extimating_unit_RST1_int), .A2(extimating_unit_RST_BLKy_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_count_RST) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_U5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_y0_int_0__5_), .B(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_block_num[1]), .Z(extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_n4)
         );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_U4 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_y0_int_0__4_), .B(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_block_num[0]), .Z(extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_n3)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurRep_U2 ( 
        .A(extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurRep_n1) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurRep_U3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_y0_int_0__3_), .B(
        extimating_unit_CE_REPy_int), .Z(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurRep_n3) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurRep_tmp_reg ( 
        .D(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurRep_n3), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurRep_n1), .Q(extimating_unit_Pixel_Retrieval_Unit_y0_int_0__3_) );
  XNOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_U6 ( 
        .A(extimating_unit_CE_BLKy_int), .B(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_0__4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n8) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_U5 ( 
        .A1(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_count_RST), .A2(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n8), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n6) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_U4 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_y0_int_0__4_), .A2(
        extimating_unit_CE_BLKy_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n9) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_U3 ( 
        .A1(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_count_RST), .A2(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n7) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_U7 ( 
        .A(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n9), .B(extimating_unit_Pixel_Retrieval_Unit_y0_int_0__5_), .Z(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n10) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_count_tmp_reg_1_ ( 
        .D(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n7), .CK(clk), .Q(extimating_unit_Pixel_Retrieval_Unit_y0_int_0__5_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_count_tmp_reg_0_ ( 
        .D(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_CurBlock_n6), .CK(clk), .Q(extimating_unit_Pixel_Retrieval_Unit_y0_int_0__4_) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_encoder_U1 ( 
        .A(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_block_num[1]), .B(extimating_unit_Pixel_Retrieval_Unit_CurCU_h_short_0_), .Z(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_y_block_num[0]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_U3 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_0__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_1__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_0__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_1__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_0__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_1__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_0__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_1__5_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_Q_int_reg_0_ ( .D(
        1'b0), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_1__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_Q_int_reg_1_ ( .D(
        1'b0), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_1__1_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_U3 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_Q_int_reg_0_ ( .D(
        1'b0), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_1__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_Q_int_reg_1_ ( .D(
        1'b0), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_1__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_0__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_1__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_0__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_1__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_0__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_1__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_0__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_1__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_1__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_2__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_1__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_2__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_1__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_2__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_1__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_2__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_1__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_2__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_1__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_2__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_1__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_2__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_1__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_2__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_1__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_2__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_1__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_2__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_1__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_2__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_1__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_2__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_2__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_3__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_2__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_3__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_2__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_3__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_2__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_3__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_2__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_3__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_2__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_3__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_2__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_3__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_2__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_3__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_2__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_3__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_2__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_3__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_2__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_3__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_2__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_3__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_3__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_3__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_3__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_3__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_3__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_3__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_4_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_3__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_3__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_3__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_3__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_3__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_3__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_4_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_5__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_5__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_5__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_5__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_5__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_5_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_5__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_5__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_5__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_5__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_5__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_5__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_5_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_5__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_5__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_6__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_5__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_6__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_5__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_6__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_5__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_6__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_5__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_6__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_5__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_6_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_6__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_5__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_6__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_5__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_6__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_5__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_6__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_5__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_6__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_5__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_6__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_5__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_6_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_6__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_6__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_7__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_6__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_7__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_6__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_7__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_6__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_7__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_6__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_7__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_6__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_7_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_7__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_6__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_7__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_6__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_7__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_6__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_7__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_6__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_7__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_6__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_7__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_6__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_7_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_7__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_7__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_8__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_7__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_8__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_7__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_8__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_7__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_8__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_7__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_8__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_7__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_8_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_8__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_7__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_8__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_7__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_8__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_7__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_8__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_7__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_8__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_7__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_8__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_7__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_8_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_8__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_8__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_9__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_8__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_9__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_8__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_9__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_8__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_9__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_8__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_9__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_8__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_9_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_9__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_8__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_9__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_8__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_9__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_8__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_9__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_8__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_9__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_8__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_9__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_8__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_9_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_9__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_9__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_10__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_9__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_10__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_9__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_10__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_9__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_10__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_9__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_10__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_9__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_10_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_10__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_9__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_10__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_9__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_10__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_9__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_10__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_9__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_10__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_9__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_10__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_9__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_10_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_10__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_10__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_11__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_10__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_11__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_10__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_11__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_10__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_11__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_10__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_11__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_10__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_11_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x0_int_11__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_10__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_11__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_10__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_11__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_10__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_11__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_10__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_11__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_10__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_11__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_10__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_11_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_11__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_11__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x_0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_11__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x_1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_11__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x_2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_11__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x_3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_11__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x_4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x0_int_11__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_X0_REG_N_X_12_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_x_5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_11__0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__0_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_11__1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_11__2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_11__3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_11__4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y0_int_11__5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_Y0_REG_N_X_12_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y0_int_12__5_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U14 ( .A(
        extimating_unit_MV0_out_int[10]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n2) );
  XNOR2_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n12), .B(
        extimating_unit_MV1_out_int[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[0]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U12 ( .A(
        extimating_unit_MV1_out_int[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n1) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U11 ( .A1(
        extimating_unit_MV0_out_int[0]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[1]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U10 ( .A(
        extimating_unit_MV0_out_int[1]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n11) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U9 ( .A(
        extimating_unit_MV0_out_int[9]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n3) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U8 ( .A(
        extimating_unit_MV0_out_int[8]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n4) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U7 ( .A(
        extimating_unit_MV0_out_int[7]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U6 ( .A(
        extimating_unit_MV0_out_int[6]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U5 ( .A(
        extimating_unit_MV0_out_int[5]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U4 ( .A(
        extimating_unit_MV0_out_int[4]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U3 ( .A(
        extimating_unit_MV0_out_int[3]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n9) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U2 ( .A(
        extimating_unit_MV0_out_int[2]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n10) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U1 ( .A(
        extimating_unit_MV0_out_int[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n12) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U2_1 ( .A(
        extimating_unit_MV1_out_int[1]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n11), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[1]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[2]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[1]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U2_2 ( .A(
        extimating_unit_MV1_out_int[2]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n10), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[2]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[3]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[2]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U2_3 ( .A(
        extimating_unit_MV1_out_int[3]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n9), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[3]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[4]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[3]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U2_4 ( .A(
        extimating_unit_MV1_out_int[4]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n8), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[4]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[5]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[4]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U2_5 ( .A(
        extimating_unit_MV1_out_int[5]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n7), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[5]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[6]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[5]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U2_6 ( .A(
        extimating_unit_MV1_out_int[6]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n6), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[6]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[7]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[6]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U2_7 ( .A(
        extimating_unit_MV1_out_int[7]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n5), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[7]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[8]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[7]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U2_8 ( .A(
        extimating_unit_MV1_out_int[8]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n4), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[8]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[9]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[8]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U2_9 ( .A(
        extimating_unit_MV1_out_int[9]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n3), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[9]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[10]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[9]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U2_10 ( .A(
        extimating_unit_MV1_out_int[10]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n2), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[10]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[11]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[10]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_U2_11 ( .A(
        extimating_unit_MV1_out_int[10]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_n2), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_0_sub_19_carry[11]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[11]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_U3 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[0]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[0]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[1]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[2]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[3]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[4]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[5]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[6]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[7]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[8]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[9]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[10]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[11]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_0_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[11]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_0_U3 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_0_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_0_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_CurCU_w_short_0_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_0_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[0]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_0_Q_int_reg_1_ ( 
        .D(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_block_num[1]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_0_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[1]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U14 ( .A(
        extimating_unit_MV0_out_int[21]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n2) );
  XNOR2_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n12), .B(
        extimating_unit_MV1_out_int[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[12]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U12 ( .A(
        extimating_unit_MV1_out_int[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n1) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U11 ( .A1(
        extimating_unit_MV0_out_int[11]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[1]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U10 ( .A(
        extimating_unit_MV0_out_int[12]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n11) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U9 ( .A(
        extimating_unit_MV0_out_int[20]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n3) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U8 ( .A(
        extimating_unit_MV0_out_int[19]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n4) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U7 ( .A(
        extimating_unit_MV0_out_int[18]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U6 ( .A(
        extimating_unit_MV0_out_int[17]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U5 ( .A(
        extimating_unit_MV0_out_int[16]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U4 ( .A(
        extimating_unit_MV0_out_int[15]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U3 ( .A(
        extimating_unit_MV0_out_int[14]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n9) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U2 ( .A(
        extimating_unit_MV0_out_int[13]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n10) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U1 ( .A(
        extimating_unit_MV0_out_int[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n12) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U2_1 ( .A(
        extimating_unit_MV1_out_int[12]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n11), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[1]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[2]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[13]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U2_2 ( .A(
        extimating_unit_MV1_out_int[13]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n10), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[2]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[3]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[14]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U2_3 ( .A(
        extimating_unit_MV1_out_int[14]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n9), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[3]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[4]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[15]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U2_4 ( .A(
        extimating_unit_MV1_out_int[15]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n8), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[4]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[5]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[16]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U2_5 ( .A(
        extimating_unit_MV1_out_int[16]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n7), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[5]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[6]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[17]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U2_6 ( .A(
        extimating_unit_MV1_out_int[17]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n6), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[6]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[7]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[18]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U2_7 ( .A(
        extimating_unit_MV1_out_int[18]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n5), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[7]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[8]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[19]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U2_8 ( .A(
        extimating_unit_MV1_out_int[19]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n4), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[8]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[9]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[20]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U2_9 ( .A(
        extimating_unit_MV1_out_int[20]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n3), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[9]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[10]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[21]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U2_10 ( .A(
        extimating_unit_MV1_out_int[21]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n2), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[10]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[11]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[22]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_U2_11 ( .A(
        extimating_unit_MV1_out_int[21]), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_n2), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_1_sub_19_carry[11]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[23]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_U3 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[12]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[12]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[13]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[13]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[14]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[14]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[15]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[15]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[16]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[16]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[17]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[17]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[18]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[18]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[19]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[19]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[20]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[20]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[21]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[21]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[22]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[22]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[23]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[23]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_1_U3 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_1_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_1_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_CurCU_w_short_0_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_1_Q_int_reg_1_ ( 
        .D(
        extimating_unit_Pixel_Retrieval_Unit_firstPelPos_calc_firstPelPos_x_block_num[1]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_1_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[3]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U14 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__9_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n3) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__8_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n4) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U12 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__7_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__5_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__3_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n9) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__2_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n10) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U6 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__10_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n2) );
  XNOR2_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n12), .B(
        extimating_unit_Pixel_Retrieval_Unit_n128), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[24]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n128), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n1) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n12) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U2 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__0_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[1]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U1 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_2__1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n11) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U2_1 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n127), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n11), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[1]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[2]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[25]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U2_2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n126), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n10), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[2]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[3]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[26]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U2_3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n125), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n9), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[3]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[4]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[27]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U2_4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n124), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n8), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[4]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[5]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[28]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U2_5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n123), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n7), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[5]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[6]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[29]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U2_6 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n122), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n6), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[6]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[7]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[30]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U2_7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n121), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n5), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[7]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[8]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[31]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U2_8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n120), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n4), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[8]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[9]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[32]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U2_9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n119), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n3), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[9]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[10]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[33]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U2_10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n118), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n2), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[10]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[11]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[34]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_U2_11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n118), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_n2), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_2_sub_19_carry[11]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[35]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_U3 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[24]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[24]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[25]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[25]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[26]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[26]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[27]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[27]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[28]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[28]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[29]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[29]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[30]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[30]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[31]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[31]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[32]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[32]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[33]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[33]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[34]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[34]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[35]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[35]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_2_U3 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_2_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_2_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_n130), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_2_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_n129), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[5]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U14 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__9_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n3) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__8_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n4) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U12 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__7_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__5_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__3_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n9) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__2_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n10) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U6 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__10_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n2) );
  XNOR2_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n12), .B(
        extimating_unit_Pixel_Retrieval_Unit_n71), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[36]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n71), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n1) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U3 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__0_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[1]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n11) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U1 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_neg_in_3__0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n12) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U2_1 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n70), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n11), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[1]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[2]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[37]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U2_2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n69), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n10), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[2]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[3]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[38]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U2_3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n68), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n9), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[3]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[4]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[39]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U2_4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n67), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n8), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[4]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[5]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[40]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U2_5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n66), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n7), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[5]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[6]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[41]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U2_6 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n65), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n6), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[6]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[7]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[42]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U2_7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n64), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n5), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[7]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[8]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[43]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U2_8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n63), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n4), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[8]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[9]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[44]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U2_9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n62), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n3), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[9]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[10]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[45]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U2_10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n61), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n2), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[10]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[11]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[46]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_U2_11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n61), .B(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_n2), .CI(
        extimating_unit_Pixel_Retrieval_Unit_SUB1_x_3_sub_19_carry[11]), .S(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[47]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_U3 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[36]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[36]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[37]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[37]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[38]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[38]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[39]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[39]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[40]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[40]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[41]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[41]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[42]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[42]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[43]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[43]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[44]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[44]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[45]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[45]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[46]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[46]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_sub1_out_tmp[47]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_SUB_OUT_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[47]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_3_U3 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_3_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_3_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_n130), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_3_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_n129), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp_x_3_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[7]) );
  OR2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_U1 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[0]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[1]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_en1) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U40 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U39 ( 
        .A(1'b1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n16) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U38 ( 
        .A1(1'b1), .A2(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[11]), 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n16), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[11]), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n52)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U37 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n52), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n2)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U36 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[10]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U35 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[9]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U34 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[8]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U33 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[7]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U32 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[6]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n9) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U31 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[5]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n10) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U30 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[4]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n11) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U29 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[3]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n12) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U28 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[2]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n13) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U27 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[1]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n14) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U26 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_en1), .A2(1'b1), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U25 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n4) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U24 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[10]), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n53)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U23 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n5), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n4), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n53), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n41)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U22 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[9]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n54)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U21 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n6), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n5), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n54), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n42)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U20 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n55)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U19 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n7), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n6), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n55), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n43)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U18 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[7]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n56)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U17 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n8), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n7), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n56), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n44)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U16 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[6]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n57)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U15 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n9), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n8), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n57), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n45)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U14 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[5]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n58)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U13 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n10), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n9), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n58), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n46)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U12 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n59)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U11 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n11), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n10), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n59), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n47)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U10 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[3]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n60)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U9 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n12), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n11), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n60), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n48)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U8 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n61)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U7 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n13), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n12), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n61), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n49)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U6 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[1]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n62)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U5 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n14), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n13), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n62), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n50)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n15) );
  OAI222_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U3 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n65), 
        .A2(1'b1), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n15), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n64), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n14), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n51)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_U2 ( 
        .A1(1'b1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n64)
         );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_SH_out_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n51), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[0]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n65) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_SH_out_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n50), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_SH_out_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n49), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_SH_out_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n48), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_SH_out_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n47), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_SH_out_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n46), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_SH_out_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n45), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_SH_out_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n44), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_SH_out_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n43), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_SH_out_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n42), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_SH_out_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n41), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_SH_out_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n2), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[11]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_en2_gen_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_en2_gen_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_en2_gen_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[1]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_en2_gen_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_en2) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U40 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U39 ( 
        .A(1'b1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n16) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U38 ( 
        .A1(1'b1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[11]), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n16), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n52) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U37 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n52), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n4)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U36 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[10]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U35 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[9]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U34 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[8]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U33 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[7]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U32 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[6]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n9) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U31 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[5]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n10) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U30 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[4]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n11) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U29 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[3]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n12) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U28 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[2]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n13) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U27 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[1]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n14) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U26 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n2) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U25 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[10]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n53)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U24 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n5), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n2), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n53), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n41)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U23 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[9]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n54)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U22 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n6), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n5), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n54), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n42)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U21 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n55)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U20 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n7), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n6), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n55), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n43)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U19 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[7]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n56)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U18 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n8), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n7), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n56), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n44)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U17 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[6]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n57)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U16 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n9), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n8), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n57), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n45)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U15 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[5]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n58)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U14 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n10), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n9), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n58), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n46)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U13 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n59)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U12 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n11), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n10), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n59), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n47)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U11 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[3]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n60)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U10 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n12), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n11), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n60), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n48)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U9 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n61)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U8 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n13), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n12), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n61), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n49)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U7 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[1]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n62)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U6 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n14), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n13), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n62), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n50)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_in_int[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n15) );
  OAI222_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U4 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n65), 
        .A2(1'b1), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n15), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n64), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n14), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n51)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U3 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_SH_en2), .A2(1'b1), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_U2 ( 
        .A1(1'b1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n64)
         );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_SH_out_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n51), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[0]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n65) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_SH_out_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n50), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_SH_out_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n49), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_SH_out_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n48), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_SH_out_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n47), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_SH_out_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n46), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_SH_out_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n45), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_SH_out_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n44), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_SH_out_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n43), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_SH_out_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n42), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_SH_out_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n41), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_SH_out_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n4), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_0_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[11]) );
  OR2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_U1 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[3]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_en1) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U40 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U39 ( 
        .A(1'b1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n16) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U38 ( 
        .A1(1'b1), .A2(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[23]), 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n16), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[11]), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n52)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U37 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n52), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n2)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U36 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[22]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U35 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[21]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U34 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[20]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U33 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[19]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U32 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[18]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n9) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U31 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[17]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n10) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U30 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[16]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n11) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U29 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[15]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n12) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U28 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[14]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n13) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U27 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[13]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n14) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U26 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_en1), .A2(1'b1), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U25 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[23]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n4) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U24 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[10]), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n53)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U23 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n5), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n4), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n53), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n41)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U22 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[9]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n54)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U21 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n6), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n5), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n54), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n42)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U20 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n55)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U19 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n7), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n6), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n55), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n43)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U18 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[7]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n56)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U17 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n8), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n7), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n56), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n44)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U16 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[6]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n57)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U15 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n9), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n8), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n57), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n45)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U14 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[5]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n58)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U13 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n10), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n9), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n58), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n46)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U12 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n59)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U11 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n11), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n10), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n59), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n47)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U10 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[3]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n60)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U9 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n12), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n11), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n60), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n48)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U8 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n61)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U7 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n13), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n12), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n61), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n49)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U6 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[1]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n62)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U5 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n14), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n13), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n62), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n50)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[12]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n15) );
  OAI222_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U3 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n65), 
        .A2(1'b1), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n15), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n64), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n14), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n51)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_U2 ( 
        .A1(1'b1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n64)
         );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_SH_out_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n51), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[0]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n65) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_SH_out_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n50), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_SH_out_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n49), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_SH_out_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n48), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_SH_out_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n47), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_SH_out_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n46), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_SH_out_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n45), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_SH_out_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n44), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_SH_out_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n43), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_SH_out_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n42), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_SH_out_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n41), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_SH_out_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n2), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[11]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_en2_gen_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_en2_gen_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_en2_gen_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[3]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_en2_gen_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_en2) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U40 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U39 ( 
        .A(1'b1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n16) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U38 ( 
        .A1(1'b1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[11]), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n16), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[23]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n52) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U37 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n52), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n4)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U36 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[10]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U35 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[9]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U34 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[8]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U33 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[7]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U32 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[6]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n9) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U31 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[5]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n10) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U30 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[4]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n11) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U29 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[3]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n12) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U28 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[2]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n13) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U27 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[1]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n14) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U26 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n2) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U25 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[22]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n53)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U24 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n5), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n2), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n53), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n41)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U23 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[21]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n54)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U22 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n6), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n5), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n54), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n42)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U21 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[20]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n55)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U20 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n7), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n6), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n55), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n43)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U19 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[19]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n56)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U18 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n8), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n7), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n56), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n44)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U17 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[18]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n57)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U16 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n9), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n8), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n57), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n45)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U15 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[17]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n58)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U14 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n10), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n9), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n58), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n46)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U13 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[16]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n59)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U12 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n11), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n10), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n59), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n47)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U11 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[15]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n60)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U10 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n12), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n11), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n60), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n48)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U9 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[14]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n61)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U8 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n13), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n12), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n61), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n49)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U7 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[13]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n62)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U6 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n14), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n13), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n62), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n50)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_in_int[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n15) );
  OAI222_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U4 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n65), 
        .A2(1'b1), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n15), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n64), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n14), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n51)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U3 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_SH_en2), .A2(1'b1), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_U2 ( 
        .A1(1'b1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n64)
         );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_SH_out_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n51), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[12]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n65) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_SH_out_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n50), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[13]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_SH_out_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n49), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[14]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_SH_out_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n48), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[15]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_SH_out_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n47), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[16]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_SH_out_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n46), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[17]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_SH_out_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n45), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[18]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_SH_out_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n44), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[19]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_SH_out_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n43), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[20]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_SH_out_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n42), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[21]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_SH_out_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n41), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[22]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_SH_out_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n4), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_1_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[23]) );
  OR2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_U1 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[5]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_en1) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U40 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U39 ( 
        .A(1'b1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n16) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U38 ( 
        .A1(1'b1), .A2(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[35]), 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n16), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[11]), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n52)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U37 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n52), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n2)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U36 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[34]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U35 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[33]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U34 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[32]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U33 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[31]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U32 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[30]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n9) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U31 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[29]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n10) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U30 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[28]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n11) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U29 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[27]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n12) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U28 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[26]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n13) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U27 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[25]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n14) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U26 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_en1), .A2(1'b1), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U25 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[35]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n4) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U24 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[10]), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n53)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U23 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n5), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n4), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n53), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n41)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U22 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[9]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n54)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U21 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n6), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n5), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n54), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n42)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U20 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n55)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U19 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n7), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n6), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n55), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n43)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U18 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[7]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n56)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U17 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n8), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n7), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n56), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n44)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U16 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[6]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n57)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U15 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n9), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n8), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n57), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n45)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U14 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[5]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n58)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U13 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n10), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n9), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n58), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n46)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U12 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n59)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U11 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n11), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n10), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n59), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n47)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U10 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[3]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n60)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U9 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n12), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n11), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n60), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n48)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U8 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n61)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U7 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n13), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n12), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n61), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n49)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U6 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[1]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n62)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U5 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n14), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n13), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n62), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n50)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[24]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n15) );
  OAI222_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U3 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n65), 
        .A2(1'b1), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n15), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n64), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n14), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n51)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_U2 ( 
        .A1(1'b1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n64)
         );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_SH_out_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n51), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[0]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n65) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_SH_out_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n50), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_SH_out_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n49), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_SH_out_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n48), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_SH_out_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n47), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_SH_out_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n46), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_SH_out_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n45), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_SH_out_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n44), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_SH_out_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n43), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_SH_out_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n42), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_SH_out_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n41), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_SH_out_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n2), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[11]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_en2_gen_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_en2_gen_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_en2_gen_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[5]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_en2_gen_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_en2) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U40 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U39 ( 
        .A(1'b1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n16) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U38 ( 
        .A1(1'b1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[11]), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n16), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__11_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n52) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U37 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n52), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n4)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U36 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[10]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U35 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[9]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U34 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[8]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U33 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[7]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U32 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[6]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n9) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U31 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[5]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n10) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U30 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[4]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n11) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U29 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[3]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n12) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U28 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[2]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n13) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U27 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[1]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n14) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U26 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n2) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U25 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__10_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n53)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U24 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n5), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n2), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n53), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n41)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U23 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__9_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n54)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U22 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n6), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n5), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n54), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n42)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U21 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__8_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n55)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U20 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n7), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n6), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n55), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n43)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U19 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__7_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n56)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U18 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n8), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n7), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n56), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n44)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U17 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n57)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U16 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n9), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n8), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n57), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n45)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U15 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__5_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n58)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U14 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n10), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n9), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n58), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n46)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U13 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__4_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n59)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U12 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n11), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n10), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n59), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n47)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U11 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__3_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n60)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U10 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n12), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n11), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n60), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n48)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U9 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__2_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n61)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U8 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n13), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n12), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n61), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n49)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U7 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__1_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n62)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U6 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n14), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n13), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n62), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n50)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_in_int[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n15) );
  OAI222_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U4 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n65), 
        .A2(1'b1), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n15), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n64), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n14), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n51)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U3 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_SH_en2), .A2(1'b1), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_U2 ( 
        .A1(1'b1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n64)
         );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_SH_out_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n51), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__0_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n65) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_SH_out_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n50), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__1_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_SH_out_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n49), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__2_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_SH_out_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n48), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__3_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_SH_out_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n47), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__4_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_SH_out_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n46), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__5_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_SH_out_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n45), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__6_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_SH_out_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n44), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__7_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_SH_out_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n43), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__8_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_SH_out_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n42), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__9_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_SH_out_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n41), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__10_) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_SH_out_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n4), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_2_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_tmp_2__11_) );
  OR2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_U1 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[6]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[7]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_en1) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U40 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U39 ( 
        .A(1'b1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n16) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U38 ( 
        .A1(1'b1), .A2(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[47]), 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n16), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[11]), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n52)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U37 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n52), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n2)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U36 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[46]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U35 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[45]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U34 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[44]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U33 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[43]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U32 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[42]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n9) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U31 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[41]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n10) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U30 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[40]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n11) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U29 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[39]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n12) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U28 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[38]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n13) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U27 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[37]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n14) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U26 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_en1), .A2(1'b1), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U25 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[47]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n4) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U24 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[10]), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n53)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U23 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n5), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n4), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n53), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n41)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U22 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[9]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n54)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U21 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n6), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n5), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n54), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n42)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U20 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n55)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U19 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n7), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n6), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n55), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n43)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U18 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[7]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n56)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U17 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n8), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n7), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n56), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n44)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U16 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[6]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n57)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U15 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n9), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n8), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n57), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n45)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U14 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[5]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n58)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U13 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n10), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n9), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n58), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n46)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U12 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n59)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U11 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n11), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n10), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n59), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n47)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U10 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[3]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n60)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U9 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n12), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n11), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n60), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n48)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U8 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n61)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U7 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n13), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n12), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n61), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n49)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U6 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[1]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n62)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U5 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n14), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n13), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n62), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n50)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_sub1_out_samp[36]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n15) );
  OAI222_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U3 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n65), 
        .A2(1'b1), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n15), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n64), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n14), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n51)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_U2 ( 
        .A1(1'b1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n64)
         );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_SH_out_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n51), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[0]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n65) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_SH_out_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n50), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_SH_out_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n49), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_SH_out_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n48), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_SH_out_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n47), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_SH_out_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n46), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_SH_out_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n45), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_SH_out_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n44), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_SH_out_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n43), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_SH_out_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n42), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_SH_out_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n41), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_SH_out_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n2), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_first_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[11]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_en2_gen_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_en2_gen_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_en2_gen_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_cmd_samp[7]), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_en2_gen_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_en2) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U40 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U39 ( 
        .A(1'b1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n16) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U38 ( 
        .A1(1'b1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[11]), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n16), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[47]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n52) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U37 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n52), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n4)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U36 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[10]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U35 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[9]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U34 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[8]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U33 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[7]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U32 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[6]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n9) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U31 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[5]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n10) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U30 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[4]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n11) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U29 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[3]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n12) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U28 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[2]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n13) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U27 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[1]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n14) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U26 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n2) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U25 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[46]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n53)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U24 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n5), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n2), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n53), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n41)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U23 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[45]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n54)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U22 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n6), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n5), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n54), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n42)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U21 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[44]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n55)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U20 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n7), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n6), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n55), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n43)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U19 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[43]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n56)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U18 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n8), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n7), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n56), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n44)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U17 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[42]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n57)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U16 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n9), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n8), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n57), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n45)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U15 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[41]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n58)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U14 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n10), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n9), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n58), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n46)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U13 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[40]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n59)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U12 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n11), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n10), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n59), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n47)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U11 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[39]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n60)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U10 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n12), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n11), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n60), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n48)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U9 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[38]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n61)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U8 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n13), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n12), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n61), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n49)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U7 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[37]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n62)
         );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U6 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n64), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n14), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n13), 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n62), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n50)
         );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_in_int[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n15) );
  OAI222_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U4 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n65), 
        .A2(1'b1), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n15), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n64), 
        .C1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n14), 
        .C2(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n51)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U3 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_SH_en2), .A2(1'b1), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_U2 ( 
        .A1(1'b1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n64)
         );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_SH_out_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n51), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[36]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n65) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_SH_out_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n50), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[37]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_SH_out_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n49), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[38]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_SH_out_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n48), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[39]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_SH_out_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n47), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[40]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_SH_out_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n46), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[41]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_SH_out_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n45), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[42]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_SH_out_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n44), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[43]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_SH_out_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n43), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[44]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_SH_out_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n42), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[45]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_SH_out_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n41), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[46]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_SH_out_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n4), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_X_3_second_shifter_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[47]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U28 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U27 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[10]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n11) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U26 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n23), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n35) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U25 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[9]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n10) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U24 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n22), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n34) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U23 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n9) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U22 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n21), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n9), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n33) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U21 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[7]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n8) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U20 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n20), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n8), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n32) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U19 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[6]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n7) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U18 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n19), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n7), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n31) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U17 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[5]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n6) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U16 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n18), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n6), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n30) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U15 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n5) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U14 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n17), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n5), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n29) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U13 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[3]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n4) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U12 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n16), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n4), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n28) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U11 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n3) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U10 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n15), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n3), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n27) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U9 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[1]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n2) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U8 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n14), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n2), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n26) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U7 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[11]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n12) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U6 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n24), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n37) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U5 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n1) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U4 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n13), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n25) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U3 ( .A(LE_ab), .Z(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n39) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_U2 ( .A(LE_ab), .Z(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n38) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n37), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[11]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n24) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n26), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[1]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n14) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n27), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[2]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n15) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n28), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[3]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n16) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n29), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[4]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n17) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n30), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[5]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n18) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_Q_int_reg_6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n31), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[6]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n19) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_Q_int_reg_7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n32), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[7]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n20) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_Q_int_reg_8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n33), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[8]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n21) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_Q_int_reg_9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n34), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[9]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n22) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n35), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[10]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n23) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n25), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[0]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_0_n13) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U28 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U27 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[22]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n65) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U26 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n53), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n65), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n41) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U25 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[21]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n66) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U24 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n54), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n66), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n42) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U23 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[20]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n67) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U22 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n55), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n67), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n43) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U21 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[19]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n68) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U20 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n56), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n68), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n44) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U19 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[18]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n69) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U18 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n57), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n69), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n45) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U17 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[17]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n70) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U16 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n58), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n70), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n46) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U15 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[16]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n71) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U14 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n59), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n71), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n47) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U13 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[15]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n72) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U12 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n60), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n72), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n48) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U11 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[14]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n73) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U10 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n61), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n73), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n49) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U9 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[13]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n74) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U8 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n62), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n74), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n50) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U7 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[12]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n75) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U6 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n63), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n51) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U5 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[23]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n64) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U4 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n52), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n40) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U3 ( .A(LE_ab), .Z(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n39) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_U2 ( .A(LE_ab), .Z(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n38) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n51), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[12]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n63) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n50), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[13]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n62) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n49), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[14]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n61) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n48), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[15]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n60) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n47), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[16]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n59) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n46), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[17]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n58) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_Q_int_reg_6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n45), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[18]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n57) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_Q_int_reg_7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n44), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[19]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n56) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_Q_int_reg_8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n43), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[20]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n55) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_Q_int_reg_9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n42), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[21]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n54) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n41), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[22]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n53) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n40), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[23]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_1_n52) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U28 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U27 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[33]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n66) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U26 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n54), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n66), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n42) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U25 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[32]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n67) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U24 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n55), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n67), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n43) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U23 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[31]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n68) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U22 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n56), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n68), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n44) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U21 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[30]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n69) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U20 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n57), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n69), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n45) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U19 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[29]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n70) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U18 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n58), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n70), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n46) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U17 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[28]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n71) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U16 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n59), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n71), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n47) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U15 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[27]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n72) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U14 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n60), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n72), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n48) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U13 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[26]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n73) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U12 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n61), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n73), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n49) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U11 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[25]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n74) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U10 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n62), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n74), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n50) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U9 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[24]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n75) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U8 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n63), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n51) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U7 ( .A(LE_ab), .Z(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U6 ( .A(LE_ab), .Z(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U5 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[34]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n65) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U4 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n53), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n65), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n41) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U3 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[35]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n64) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_U2 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n52), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n38), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n40) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n51), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[24]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n63) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n50), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[25]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n62) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n49), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[26]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n61) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n48), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[27]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n60) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n47), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[28]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n59) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n46), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[29]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n58) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_Q_int_reg_6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n45), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[30]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n57) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_Q_int_reg_7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n44), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[31]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n56) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_Q_int_reg_8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n43), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[32]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n55) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_Q_int_reg_9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n42), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[33]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n54) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n41), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[34]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n53) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n40), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[35]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_2_n52) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U28 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U27 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[46]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n65) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U26 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n53), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n65), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n41) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U25 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[45]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n66) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U24 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n54), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n66), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n42) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U23 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[44]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n67) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U22 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n55), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n67), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n43) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U21 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[43]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n68) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U20 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n56), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n68), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n44) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U19 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[42]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n69) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U18 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n57), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n69), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n45) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U17 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[41]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n70) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U16 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n58), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n70), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n46) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U15 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[40]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n71) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U14 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n59), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n71), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n47) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U13 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[39]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n72) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U12 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n60), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n72), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n48) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U11 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[38]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n73) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U10 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n61), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n73), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n49) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U9 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[37]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n74) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U8 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n62), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n74), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n50) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U7 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[47]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n64) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U6 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n52), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n40) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U5 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39), .A2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out[36]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n75) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U4 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n63), .B2(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39), .A(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n51) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U3 ( .A(LE_ab), .Z(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n39) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_U2 ( .A(LE_ab), .Z(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n38) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n51), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[36]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n63) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n50), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[37]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n62) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n49), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[38]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n61) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n48), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[39]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n60) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n47), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[40]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n59) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n46), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[41]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n58) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_Q_int_reg_6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n45), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[42]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n57) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_Q_int_reg_7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n44), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[43]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n56) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_Q_int_reg_8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n43), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[44]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n55) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_Q_int_reg_9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n42), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[45]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n54) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n41), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[46]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n53) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n40), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[47]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_a12b12_REG_3_n52) );
  NOR3_X4 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U103 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_int_LE), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_), .A3(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n86), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U102 ( .A1(1'b0), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op2_int_6_) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U101 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_11_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_5_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n80) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U100 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n80), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n27) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U99 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_10_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_4_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n81) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U98 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n81), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n28) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U97 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_9_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_3_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n82) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U96 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n82), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n29) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U95 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_8_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_2_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n83) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U94 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n83), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n30) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U93 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_7_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_1_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n84) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U92 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n84), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n31) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U91 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_0_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n85) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U90 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n85), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n32) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U89 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_11_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_5_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n73) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U88 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n73), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n10) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U87 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_10_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n75) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U86 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n12) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U85 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_9_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_3_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n76) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U84 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n76), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n14) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U83 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_8_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_2_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n77) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U82 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n77), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n16) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U81 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_7_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n78) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U80 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n78), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n18) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U79 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_6_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n79) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U78 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n79), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n20) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U77 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__1_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n46) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U76 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n46), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n25) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U75 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__0_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n47) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U74 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n47), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n26) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U73 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__3_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n44) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U72 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n44), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n23) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U71 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_25_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n56), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_N35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n54) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U70 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n54), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n1) );
  AOI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U69 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n41), .B2(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__5_), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n42) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U68 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n42), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n21) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U67 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__4_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n43) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U66 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n43), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n22) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U65 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__2_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n45) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U64 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n45), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n24) );
  AOI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U63 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n40), .B2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[5]), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op1_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n48) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U62 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n48), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n34) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U61 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n40), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[10]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n49) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U60 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n49), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n35) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U59 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n40), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[8]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n51) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U58 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n51), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n37) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U57 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[1]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n40), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[7]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n52) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U56 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n52), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n38) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U55 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[0]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n40), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[6]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n53) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U54 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n53), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n39) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U53 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[3]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n40), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[9]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n50) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U52 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n50), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n36) );
  OR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U51 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n36), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_rst_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n86) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U50 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_24_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n59) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U49 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n2), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n58), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n59), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n87) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U48 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_23_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n60) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U47 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n3), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n58), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n60), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n88) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U46 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_22_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n61) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U45 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n4), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n58), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n61), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n89) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U44 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_21_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n62) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U43 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n5), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n58), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n62), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n90) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U42 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_20_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n63) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U41 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n6), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n58), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n91) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U40 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_19_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n64) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U39 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n7), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n58), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n92) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U38 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[11]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op1_int_6_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U37 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n41) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U36 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_12_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n72) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U35 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n19) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U34 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n19), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n65), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n8), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n72), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n99) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U33 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_13_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n71) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U32 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n17) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U31 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n17), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n65), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n7), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n71), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n98) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U30 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_14_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n70) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U29 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_2_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n15) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U28 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n15), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n65), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n6), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n70), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n97) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U27 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_15_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n69) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_3_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n13) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U25 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n13), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n65), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n5), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n69), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n96) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U24 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_16_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n68) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U23 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n11) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U22 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n11), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n65), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n4), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n68), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n95) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U21 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_17_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n67) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U20 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_5_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n9) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U19 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n9), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n65), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n3), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n67), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n94) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U18 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_18_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n66) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U17 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n8), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n65), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n2), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n66), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n93) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U16 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n40) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U15 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n56), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n65) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U14 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n86), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n74) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U12 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_12_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n2) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_7_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_8_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_9_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_10_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n4) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_11_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n3) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U6 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_N35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n58) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U5 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n86), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n55), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n56) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n65), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n33) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_U3 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n56), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n57) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n32), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_0_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n31), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_1_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n30), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_2_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n29), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_3_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n28), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_4_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n27), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_5_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n20), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_6_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n18), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_7_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n16), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_8_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n14), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_9_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n12), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_10_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n10), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_11_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_19_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n92), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_19_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_20_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n91), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_20_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_21_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n90), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_21_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_22_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n89), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_22_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_23_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n88), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_23_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_24_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n87), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_24_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_25_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n1), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_25_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_18_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n93), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_18_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_17_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n94), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_17_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_16_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n95), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_16_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_15_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n96), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_15_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_14_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n97), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_14_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n98), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_13_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n99), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_12_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n2) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_U5 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n3), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n4), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_rst_0_) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_U4 ( 
        .A1(MULT1_VALID), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_count_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n5), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_1_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n3) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_count_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n7), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n4) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_U6 ( 
        .A(MULT1_VALID), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_count_int_0_), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n7) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_U3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n1), 
        .B(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n3), 
        .Z(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_ctrl_sign_gen_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n2) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[0]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[0]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[1]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[2]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[3]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[4]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[5]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[6]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[7]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[8]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[9]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[10]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[11]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[11]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[12]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[12]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_Q_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[13]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1_sampling_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[13]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_12_), 
        .B(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[0]), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_0_) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_12_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_n1) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1_1 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[1]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_13_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_n1), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[2]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_1_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1_2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[2]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_14_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[2]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[3]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_2_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1_3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[3]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_15_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[3]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[4]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_3_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1_4 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[4]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_16_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[4]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[5]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_4_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1_5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[5]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_17_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[5]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[6]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_5_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1_6 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[6]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_18_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[6]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[7]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_6_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1_7 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[7]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_19_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[7]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[8]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_7_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1_8 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[8]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_20_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[8]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[9]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_8_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1_9 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[9]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_21_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[9]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[10]), .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_9_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1_10 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[10]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_22_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[10]), .CO(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[11]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_10_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1_11 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[11]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_23_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[11]), .CO(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[12]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_11_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1_12 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[12]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_24_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[12]), .CO(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[13]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_12_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_U1_13 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add1[13]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_25_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_pp_sum_add_19_carry[13]), .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_N35) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_int_LE_FF_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_int_LE_FF_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_int_LE_FF_Q_int_reg ( 
        .D(MULT1_VALID), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_int_LE_FF_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_int_LE) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_RST_FFX_1_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_RST_FFX_1_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_RST_FFX_1_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_rst_0_), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_RST_FFX_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_rst_1_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_RST_FFX_2_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_RST_FFX_2_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_RST_FFX_2_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_rst_1_), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_RST_FFX_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_RST_FFX_2_Q) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_result_LE_FF_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_result_LE_FF_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_result_LE_FF_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_SUM_rst_0_), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_result_LE_FF_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_result_LE) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U56 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U55 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_5_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n6) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U54 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n30), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n6), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n54) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U53 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_4_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n5) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U52 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n29), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n5), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n53) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U51 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_3_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n4) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U50 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n28), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n4), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n52) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U49 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_2_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n3) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U48 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n27), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n3), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n51) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U47 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_1_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n2) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U46 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n26), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n2), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n50) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U45 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_5_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n18) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U44 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n42), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n18), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n66) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U43 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_result_LE), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n74) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U42 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_result_LE), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n72) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U41 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n19) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U40 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n43), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n19), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n67) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U39 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_4_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n17) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U38 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n41), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n17), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n65) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U37 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_3_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n16) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U36 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n40), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n64) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U35 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_2_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n15) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U34 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n39), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n15), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n63) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U33 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_1_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n14) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U32 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n38), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n14), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n62) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U31 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_0_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n13) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U30 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n37), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n13), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n61) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U29 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_11_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n12) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U28 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n36), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n12), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n60) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U27 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_10_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n11) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U26 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n35), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n11), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n59) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U25 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_9_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n10) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U24 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n34), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n10), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n58) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U23 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_8_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n9) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U22 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n33), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n9), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n57) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U21 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_7_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n8) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U20 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n32), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n8), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n56) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U19 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_6_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n7) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U18 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n31), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n7), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n55) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U17 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_int_0_), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n1) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U16 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n25), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n49) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U15 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_11_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n24) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U14 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n48), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n24), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n73) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U13 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_10_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n23) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U12 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n47), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n23), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n71) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U11 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_9_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n22) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U10 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n46), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n22), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n70) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U9 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_8_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n21) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U8 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n45), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n21), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n69) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U7 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_add_out_7_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n20) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U6 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n44), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n20), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n68) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n74), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n78) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n74), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n77) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n72), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n76) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_U2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n72), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n75) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_23_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n73), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_23_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n48) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_22_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n71), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_22_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n47) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_21_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n70), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_21_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n46) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_20_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n69), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_20_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n45) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_19_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n68), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_19_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n44) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_18_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n67), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_product_18_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n43) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_17_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n66), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[17]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n42) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_16_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n65), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[16]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n41) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_15_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n64), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[15]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n40) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_14_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n63), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[14]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n39) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n62), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[13]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n38) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n61), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[12]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n37) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n57), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[8]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n33) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n50), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[1]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n26) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n51), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[2]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n27) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n52), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[3]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n28) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n55), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[6]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n31) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n53), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[4]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n29) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n54), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[5]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n30) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n56), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[7]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n32) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n58), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[9]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n34) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n59), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[10]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n35) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n60), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[11]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n36) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n49), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[0]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_output_reg_n25) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U173 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n176), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n100) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U172 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n37), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n101) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U171 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n168), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n177), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n102) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U170 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n169), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n177), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n103) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U169 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n177), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n104) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U168 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n171), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n177), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n105) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U167 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n172), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n177), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n106) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U166 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n177), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n107) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U165 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n38), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n108) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U164 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n168), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n178), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n109) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U163 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n169), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n178), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n110) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U162 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n178), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n111) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U161 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n171), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n178), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n112) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U160 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n172), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n178), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n113) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U159 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n178), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n114) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U158 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op2_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n115) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U157 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n116) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U156 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n117) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U155 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n170), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n118) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U154 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n119) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U153 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n120) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U152 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n22), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n181) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U151 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n34), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n24), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n180) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U150 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n181), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n180), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n41) );
  XNOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U149 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n180), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n181), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n42) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U148 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op2_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op1_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n73) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U147 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n21), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n74) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U146 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n22), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n75) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U145 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n76) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U144 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n24), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n77) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U143 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n25), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n78) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U142 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n26), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n79) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U141 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n34), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n80) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U140 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n168), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n174), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n81) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U139 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n169), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n174), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n82) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U138 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n174), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n83) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U137 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n172), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n174), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n85) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U136 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n174), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n86) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U135 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n35), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n87) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U134 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n168), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n175), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n88) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U133 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n175), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n89) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U132 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n175), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n90) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U131 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n171), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n175), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n91) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U130 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n172), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n175), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n92) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U129 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n175), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n93) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U128 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_op2_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n94) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U127 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n95) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U126 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n170), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n97) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U125 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n98) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U124 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n99) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U123 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n173), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[0]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U122 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n34), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n174) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U121 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n22), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n169) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U120 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n24), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n171) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U119 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n176) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U118 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n178) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U117 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n177) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U116 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n175) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U115 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n21), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n168) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U114 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n170) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U113 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n25), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n172) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U112 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n26), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n173) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U111 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n179) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U110 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[13]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U44 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n113), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n119), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n71), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n72) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U43 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n100), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n106), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n69), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n70) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U42 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n112), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n118), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n71), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n67), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n68) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U41 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n93), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n99), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n65), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n66) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U40 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n105), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n117), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n111), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n63), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n64) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U39 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n66), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n69), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n67), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n61), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n62) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U38 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n86), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n92), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n59), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n60) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U37 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n98), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n116), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n104), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n57), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n58) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U36 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n65), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n110), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n60), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n55), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n56) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U35 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n58), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n63), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n56), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n53), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n54) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U34 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n97), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n91), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n51), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n52) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U33 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n85), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n103), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n109), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n49), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n50) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U32 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n79), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n115), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n59), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n47), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n48) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U31 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n57), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n52), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n50), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n45), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n46) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U30 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n48), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n55), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n46), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n43), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n44) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U27 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n102), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n90), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n108), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n39), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n40) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n51), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n78), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n42), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n37), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n38) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U25 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n47), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n49), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n40), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n35), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n36) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U24 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n45), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n38), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n36), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n33), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n34) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U23 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n83), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n89), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n95), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n31), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n32) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U22 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n77), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n101), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n41), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n29), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n30) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U21 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n32), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n39), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n37), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n27), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n28) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U20 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n35), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n30), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n28), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n25), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n26) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U19 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n82), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n88), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n94), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n23), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n24) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U18 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n31), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n76), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n29), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n21), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n22) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U17 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n27), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n24), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n22), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n19), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n20) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U16 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n87), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n81), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n75), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n17), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n18) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U15 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n18), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n23), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n21), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n15), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n16) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U14 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n74), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n80), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n17), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n13), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n14) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n120), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n114), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n12), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[1]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U12 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n12), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n107), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n72), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n11), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[2]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n11), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n70), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n68), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n10), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[3]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n62), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n64), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n10), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n9), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[4]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n54), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n61), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n9), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n8), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[5]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n44), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n53), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n8), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n7), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[6]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n34), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n43), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n7), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n6), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[7]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U6 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n26), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n33), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n6), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n5), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[8]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n20), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n25), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n5), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n4), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[9]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n16), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n19), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n4), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n3), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[10]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n15), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n14), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n3), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n2), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[11]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_U2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n13), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n73), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n2), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_47_n1), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_0_mult_int[12]) );
  NOR3_X4 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U103 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_int_LE), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_), .A3(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n113), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U102 ( .A1(1'b0), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op2_int_6_) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U101 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_11_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_5_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n119) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U100 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n119), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n28) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U99 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_10_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_4_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n118) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U98 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n118), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n29) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U97 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_9_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_3_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n117) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U96 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n117), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n30) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U95 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_8_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_2_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n116) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U94 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n116), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n31) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U93 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_7_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_1_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n115) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U92 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n115), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n32) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U91 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_0_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n114) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U90 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n114), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n33) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U89 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_11_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_5_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n126) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U88 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n126), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n10) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U87 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_10_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n124) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U86 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n124), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n12) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U85 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_9_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_3_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n123) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U84 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n123), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n14) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U83 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_8_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_2_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n122) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U82 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n122), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n16) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U81 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_7_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n121) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U80 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n121), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n18) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U79 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_6_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n120) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U78 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n120), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n20) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U77 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__1_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n153) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U76 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n153), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n39) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U75 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__0_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n152) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U74 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n152), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n40) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U73 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__3_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n155) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U72 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n155), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n37) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U71 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_25_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n143), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_N35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n145) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U70 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n145), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n1) );
  AOI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U69 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n41), .B2(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__5_), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n157) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U68 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n157), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n35) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U67 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__4_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n156) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U66 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n156), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n36) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U65 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_0__2_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n154) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U64 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n154), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n38) );
  AOI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U63 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n27), .B2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[17]), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op1_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n151) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U62 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n151), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n21) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U61 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[16]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[22]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n150) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U60 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n150), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n22) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U59 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[14]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[20]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n148) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U58 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n148), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n24) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U57 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[13]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[19]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n147) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U56 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n147), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n25) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U55 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[12]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[18]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n146) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U54 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n146), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n26) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U53 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[15]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[21]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n149) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U52 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n149), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n23) );
  OR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U51 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n36), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_rst_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n113) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U50 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_24_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n140) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U49 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n2), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n140), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n112) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U48 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_23_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n139) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U47 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n3), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n139), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n111) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U46 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_22_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n138) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U45 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n4), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n138), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n110) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U44 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_21_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n137) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U43 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n5), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n137), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n109) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U42 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_20_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n136) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U41 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n6), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n136), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n108) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U40 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_19_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n135) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U39 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n7), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n135), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n107) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U38 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[23]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op1_int_6_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U37 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n41) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U36 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_12_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n127) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U35 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n19) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U34 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n19), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n8), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n127), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n100) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U33 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_13_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n128) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U32 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n17) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U31 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n17), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n7), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n128), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n101) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U30 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_14_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n129) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U29 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_2_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n15) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U28 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n15), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n6), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n129), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n102) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U27 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_15_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n130) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_3_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n13) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U25 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n13), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n5), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n130), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n103) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U24 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_16_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n131) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U23 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n11) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U22 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n11), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n4), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n131), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n104) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U21 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_17_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n132) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U20 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_5_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n9) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U19 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n9), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n3), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n132), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n105) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U18 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_18_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n133) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U17 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n8), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n2), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n133), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n106) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U16 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n27) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U15 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n143), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n134) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U14 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n113), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n125) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U12 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_12_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n2) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_7_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_8_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_9_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_10_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n4) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_11_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n3) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U6 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_N35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n141) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U5 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n113), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n143) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n134), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n34) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_U3 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n143), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n27), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n142) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n33), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_0_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n32), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_1_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n31), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_2_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n30), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_3_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n29), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_4_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n28), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_5_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n20), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_6_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n18), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_7_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n16), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_8_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n14), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_9_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n12), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_10_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n10), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_11_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_19_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n107), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_19_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_20_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n108), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_20_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_21_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n109), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_21_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_22_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n110), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_22_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_23_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n111), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_23_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_24_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n112), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_24_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_25_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n1), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_25_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_18_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n106), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_18_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_17_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n105), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_17_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_16_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n104), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_16_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_15_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n103), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_15_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_14_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n102), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_14_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n101), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_13_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n100), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_12_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n2) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_U5 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n9), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n8), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_rst_0_) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_U4 ( 
        .A1(MULT1_VALID), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n10) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_U6 ( 
        .A(MULT1_VALID), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n6) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_U3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n10), 
        .B(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n9), 
        .Z(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n7) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_count_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n7), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_1_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n9) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_count_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n6), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_count_int_0_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_ctrl_sign_gen_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n2) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[0]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[0]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[1]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[2]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[3]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[4]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[5]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[6]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[7]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[8]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[9]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[10]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[11]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[11]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[12]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[12]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_Q_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[13]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1_sampling_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[13]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_12_), 
        .B(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[0]), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_0_) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_12_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_n1) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1_1 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[1]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_13_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_n1), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[2]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_1_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1_2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[2]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_14_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[2]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[3]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_2_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1_3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[3]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_15_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[3]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[4]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_3_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1_4 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[4]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_16_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[4]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[5]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_4_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1_5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[5]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_17_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[5]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[6]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_5_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1_6 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[6]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_18_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[6]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[7]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_6_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1_7 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[7]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_19_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[7]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[8]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_7_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1_8 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[8]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_20_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[8]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[9]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_8_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1_9 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[9]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_21_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[9]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[10]), .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_9_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1_10 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[10]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_22_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[10]), .CO(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[11]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_10_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1_11 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[11]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_23_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[11]), .CO(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[12]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_11_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1_12 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[12]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_24_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[12]), .CO(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[13]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_12_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_U1_13 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add1[13]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_25_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_pp_sum_add_19_carry[13]), .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_N35) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_int_LE_FF_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_int_LE_FF_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_int_LE_FF_Q_int_reg ( 
        .D(MULT1_VALID), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_int_LE_FF_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_int_LE) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_RST_FFX_1_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_RST_FFX_1_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_RST_FFX_1_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_rst_0_), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_RST_FFX_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_rst_1_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_RST_FFX_2_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_RST_FFX_2_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_RST_FFX_2_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_rst_1_), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_RST_FFX_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_RST_FFX_2_Q) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_result_LE_FF_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_result_LE_FF_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_result_LE_FF_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_SUM_rst_0_), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_result_LE_FF_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_result_LE) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U57 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U56 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U55 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_5_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n147) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U54 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n123), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n147), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n99) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U53 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_4_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n148) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U52 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n124), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n148), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n100) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U51 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_3_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n149) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U50 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n125), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n149), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n101) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U49 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_2_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n150) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U48 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n126), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n150), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n102) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U47 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_1_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n151) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U46 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n127), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n151), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n103) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U45 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_5_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n135) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U44 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n111), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n135), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n87) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U43 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_result_LE), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n74) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U42 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_result_LE), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n72) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U41 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n134) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U40 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n110), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n134), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n86) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U39 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_4_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n136) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U38 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n112), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n136), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n88) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U37 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_3_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n137) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U36 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n113), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n137), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n89) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U35 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_2_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n138) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U34 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n114), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n138), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n90) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U33 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_1_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n139) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U32 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n115), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n139), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n91) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U31 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_0_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n140) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U30 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n116), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n140), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n92) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U29 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_11_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n141) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U28 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n117), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n141), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n93) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U27 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_10_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n142) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U26 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n118), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n142), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n94) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U25 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_9_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n143) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U24 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n119), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n143), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n95) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U23 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_8_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n144) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U22 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n120), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n144), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n96) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U21 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_7_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n145) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U20 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n121), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n145), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n97) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U19 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_6_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n146) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U18 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n122), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n146), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n98) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U17 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_int_0_), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n152) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U16 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n128), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n152), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n104) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U15 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_11_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n129) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U14 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n105), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n129), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n81) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U13 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_10_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n130) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U12 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n106), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n130), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n82) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U11 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_9_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n131) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U10 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n107), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n131), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n83) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U9 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_8_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n132) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U8 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n108), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n132), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n84) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U7 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_add_out_7_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n133) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U6 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n109), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n133), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n85) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n74), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n78) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n74), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n77) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n72), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n76) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_U2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n72), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n75) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n104), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[0]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n128) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n103), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[1]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n127) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n102), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[2]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n126) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n101), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[3]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n125) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n100), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[4]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n124) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n99), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[5]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n123) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n98), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[6]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n122) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n97), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[7]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n121) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n96), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[8]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n120) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n95), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[9]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n119) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n94), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[10]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n118) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n93), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[11]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n117) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n92), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[12]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n116) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n91), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[13]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n115) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_14_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n90), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[14]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n114) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_15_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n89), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[15]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n113) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_16_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n88), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[16]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n112) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_17_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n87), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[17]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n111) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_18_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n86), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_18_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n110) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_19_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n85), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_19_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n109) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_20_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n84), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_20_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n108) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_21_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n83), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_21_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n107) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_22_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n82), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_22_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n106) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_Q_int_reg_23_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n81), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_product_23_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_output_reg_n105) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U173 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n170), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n100) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U172 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n24), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n101) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U171 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n174), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n102) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U170 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n175), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n103) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U169 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n104) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U168 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n177), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n105) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U167 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n178), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n106) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U166 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n107) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U165 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n25), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n108) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U164 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n174), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n109) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U163 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n175), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n110) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U162 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n111) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U161 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n177), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n112) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U160 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n178), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n113) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U159 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n114) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U158 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op2_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n26), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n115) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U157 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n174), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n116) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U156 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n175), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n117) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U155 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n176), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n118) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U154 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n177), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n119) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U153 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n178), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n120) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U152 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n36), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n181) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U151 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n21), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n180) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U150 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n181), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n180), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n41) );
  XNOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U149 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n180), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n181), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n42) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U148 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op2_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op1_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n73) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U147 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n74) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U146 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n75) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U145 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n76) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U144 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n77) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U143 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n78) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U142 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n79) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U141 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n21), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n80) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U140 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n174), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n81) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U139 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n175), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n82) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U138 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n83) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U137 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n178), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n85) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U136 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n86) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U135 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n22), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n87) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U134 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n174), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n88) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U133 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n169), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n175), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n89) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U132 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n90) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U131 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n177), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n91) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U130 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n178), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n92) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U129 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n93) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U128 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_op2_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n94) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U127 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n174), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n95) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U126 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n176), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n97) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U125 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n177), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n98) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U124 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n178), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n99) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U123 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n179), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[0]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U122 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n21), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n168) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U121 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n175) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U120 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n177) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U119 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n170) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U118 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n25), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n172) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U117 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n24), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n171) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U116 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n22), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n169) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U115 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n174) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U114 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n176) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U113 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n178) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U112 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n179) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U111 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_n26), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n173) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U110 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[13]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U44 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n113), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n119), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n71), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n72) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U43 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n100), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n106), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n69), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n70) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U42 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n112), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n118), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n71), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n67), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n68) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U41 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n93), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n99), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n65), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n66) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U40 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n105), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n117), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n111), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n63), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n64) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U39 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n66), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n69), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n67), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n61), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n62) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U38 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n86), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n92), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n59), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n60) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U37 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n98), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n116), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n104), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n57), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n58) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U36 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n65), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n110), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n60), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n55), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n56) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U35 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n58), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n63), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n56), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n53), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n54) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U34 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n97), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n91), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n51), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n52) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U33 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n85), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n103), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n109), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n49), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n50) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U32 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n79), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n115), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n59), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n47), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n48) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U31 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n57), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n52), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n50), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n45), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n46) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U30 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n48), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n55), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n46), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n43), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n44) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U27 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n102), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n90), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n108), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n39), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n40) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n51), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n78), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n42), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n37), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n38) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U25 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n47), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n49), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n40), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n35), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n36) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U24 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n45), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n38), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n36), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n33), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n34) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U23 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n83), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n89), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n95), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n31), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n32) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U22 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n77), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n101), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n41), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n29), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n30) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U21 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n32), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n39), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n37), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n27), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n28) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U20 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n35), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n30), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n28), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n25), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n26) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U19 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n82), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n88), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n94), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n23), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n24) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U18 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n31), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n76), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n29), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n21), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n22) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U17 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n27), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n24), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n22), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n19), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n20) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U16 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n87), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n81), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n75), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n17), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n18) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U15 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n18), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n23), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n21), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n15), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n16) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U14 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n74), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n80), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n17), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n13), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n14) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n120), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n114), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n12), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[1]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U12 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n12), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n107), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n72), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n11), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[2]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n11), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n70), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n68), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n10), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[3]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n62), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n64), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n10), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n9), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[4]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n54), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n61), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n9), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n8), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[5]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n44), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n53), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n8), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n7), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[6]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n34), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n43), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n7), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n6), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[7]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U6 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n26), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n33), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n6), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n5), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[8]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n20), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n25), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n5), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n4), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[9]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n16), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n19), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n4), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n3), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[10]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n15), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n14), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n3), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n2), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[11]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_U2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n13), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n73), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n2), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_47_n1), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_1_mult_int[12]) );
  NOR3_X4 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U103 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_int_LE), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_), .A3(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n113), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U102 ( .A1(1'b0), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op2_int_6_) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U101 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_11_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_5_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n119) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U100 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n119), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n28) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U99 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_10_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_4_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n118) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U98 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n118), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n29) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U97 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_9_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_3_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n117) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U96 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n117), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n30) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U95 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_8_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_2_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n116) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U94 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n116), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n31) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U93 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_7_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_1_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n115) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U92 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n115), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n32) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U91 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_0_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n114) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U90 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n114), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n33) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U89 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_11_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_5_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n126) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U88 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n126), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n10) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U87 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_10_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n124) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U86 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n124), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n12) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U85 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_9_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_3_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n123) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U84 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n123), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n14) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U83 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_8_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_2_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n122) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U82 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n122), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n16) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U81 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_7_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n121) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U80 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n121), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n18) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U79 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_6_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n120) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U78 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n120), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n20) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U77 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__1_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n153) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U76 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n153), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n39) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U75 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__0_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n152) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U74 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n152), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n40) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U73 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__3_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n155) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U72 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n155), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n37) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U71 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_25_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n143), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_N35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n145) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U70 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n145), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n1) );
  AOI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U69 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n41), .B2(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__5_), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n157) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U68 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n157), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n35) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U67 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__4_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n156) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U66 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n156), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n36) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U65 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__2_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n154) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U64 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n154), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n38) );
  AOI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U63 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n27), .B2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[29]), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op1_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n151) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U62 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n151), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n21) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U61 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[28]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[34]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n150) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U60 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n150), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n22) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U59 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[26]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[32]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n148) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U58 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n148), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n24) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U57 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[25]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[31]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n147) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U56 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n147), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n25) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U55 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[24]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[30]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n146) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U54 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n146), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n26) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U53 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[27]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[33]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n149) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U52 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n149), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n23) );
  OR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U51 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n36), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_rst_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n113) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U50 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_24_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n140) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U49 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n2), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n140), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n112) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U48 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_23_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n139) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U47 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n3), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n139), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n111) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U46 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_22_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n138) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U45 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n4), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n138), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n110) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U44 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_21_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n137) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U43 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n5), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n137), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n109) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U42 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_20_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n136) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U41 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n6), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n136), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n108) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U40 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_19_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n135) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U39 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n7), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n135), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n107) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U38 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[35]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op1_int_6_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U37 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n41) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U36 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_12_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n127) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U35 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n19) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U34 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n19), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n8), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n127), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n100) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U33 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_13_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n128) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U32 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n17) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U31 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n17), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n7), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n128), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n101) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U30 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_14_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n129) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U29 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_2_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n15) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U28 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n15), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n6), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n129), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n102) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U27 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_15_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n130) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_3_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n13) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U25 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n13), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n5), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n130), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n103) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U24 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_16_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n131) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U23 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n11) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U22 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n11), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n4), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n131), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n104) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U21 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_17_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n132) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U20 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_5_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n9) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U19 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n9), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n3), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n132), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n105) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U18 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_18_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n133) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U17 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n8), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n2), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n133), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n106) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U16 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n27) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U15 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n143), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n134) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U14 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n113), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n125) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U12 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_12_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n2) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_7_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_8_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_9_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_10_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n4) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_11_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n3) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U6 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_N35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n141) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U5 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n113), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n143) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n134), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n34) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_U3 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n143), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n27), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n142) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n33), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_0_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n32), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_1_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n31), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_2_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n30), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_3_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n29), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_4_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n28), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_5_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n20), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_6_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n18), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_7_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n16), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_8_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n14), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_9_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n12), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_10_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n10), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_11_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_19_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n107), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_19_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_20_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n108), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_20_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_21_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n109), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_21_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_22_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n110), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_22_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_23_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n111), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_23_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_24_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n112), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_24_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_25_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n1), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_25_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_18_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n106), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_18_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_17_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n105), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_17_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_16_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n104), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_16_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_15_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n103), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_15_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_14_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n102), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_14_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n101), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_13_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n100), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_12_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n2) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_U5 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n9), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n8), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_rst_0_) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_U4 ( 
        .A1(MULT1_VALID), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n10) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_U6 ( 
        .A(MULT1_VALID), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n6) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_U3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n10), 
        .B(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n9), 
        .Z(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n7) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_count_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n7), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_1_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n9) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_count_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n6), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_count_int_0_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_ctrl_sign_gen_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n2) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[0]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[0]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[1]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[2]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[3]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[4]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[5]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[6]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[7]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[8]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[9]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[10]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[11]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[11]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[12]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[12]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_Q_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[13]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1_sampling_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[13]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_12_), 
        .B(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[0]), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_0_) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_12_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_n1) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1_1 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[1]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_13_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_n1), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[2]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_1_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1_2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[2]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_14_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[2]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[3]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_2_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1_3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[3]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_15_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[3]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[4]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_3_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1_4 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[4]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_16_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[4]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[5]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_4_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1_5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[5]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_17_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[5]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[6]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_5_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1_6 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[6]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_18_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[6]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[7]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_6_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1_7 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[7]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_19_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[7]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[8]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_7_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1_8 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[8]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_20_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[8]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[9]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_8_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1_9 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[9]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_21_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[9]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[10]), .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_9_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1_10 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[10]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_22_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[10]), .CO(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[11]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_10_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1_11 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[11]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_23_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[11]), .CO(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[12]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_11_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1_12 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[12]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_24_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[12]), .CO(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[13]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_12_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_U1_13 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add1[13]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_25_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_pp_sum_add_19_carry[13]), .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_N35) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_int_LE_FF_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_int_LE_FF_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_int_LE_FF_Q_int_reg ( 
        .D(MULT1_VALID), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_int_LE_FF_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_int_LE) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_RST_FFX_1_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_RST_FFX_1_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_RST_FFX_1_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_rst_0_), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_RST_FFX_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_rst_1_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_RST_FFX_2_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_RST_FFX_2_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_RST_FFX_2_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_rst_1_), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_RST_FFX_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_RST_FFX_2_Q) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_result_LE_FF_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_result_LE_FF_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_result_LE_FF_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_SUM_rst_0_), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_result_LE_FF_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_result_LE) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U57 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U56 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U55 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_5_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n147) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U54 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n123), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n147), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n99) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U53 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_4_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n148) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U52 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n124), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n148), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n100) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U51 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_3_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n149) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U50 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n125), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n149), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n101) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U49 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_2_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n150) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U48 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n126), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n150), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n102) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U47 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_1_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n151) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U46 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n127), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n151), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n103) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U45 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_5_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n135) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U44 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n111), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n135), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n87) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U43 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_result_LE), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n74) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U42 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_result_LE), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n72) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U41 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n134) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U40 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n110), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n134), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n86) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U39 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_4_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n136) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U38 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n112), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n136), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n88) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U37 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_3_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n137) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U36 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n113), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n137), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n89) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U35 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_2_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n138) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U34 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n114), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n138), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n90) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U33 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_1_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n139) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U32 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n115), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n139), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n91) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U31 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_0_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n140) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U30 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n116), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n140), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n92) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U29 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_11_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n141) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U28 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n117), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n141), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n93) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U27 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_10_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n142) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U26 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n118), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n142), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n94) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U25 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_9_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n143) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U24 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n119), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n143), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n95) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U23 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_8_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n144) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U22 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n120), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n144), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n96) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U21 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_7_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n145) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U20 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n121), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n145), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n97) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U19 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_6_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n146) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U18 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n122), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n146), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n98) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U17 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_int_0_), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n152) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U16 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n128), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n152), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n104) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U15 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_11_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n129) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U14 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n105), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n129), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n81) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U13 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_10_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n130) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U12 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n106), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n130), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n82) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U11 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_9_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n131) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U10 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n107), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n131), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n83) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U9 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_8_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n132) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U8 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n108), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n132), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n84) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U7 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_add_out_7_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n133) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U6 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n109), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n133), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n85) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n74), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n78) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n74), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n77) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n72), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n76) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_U2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n72), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n75) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n104), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[0]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n128) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n103), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[1]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n127) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n102), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[2]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n126) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n101), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[3]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n125) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n100), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[4]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n124) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n99), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[5]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n123) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n98), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[6]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n122) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n97), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[7]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n121) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n96), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[8]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n120) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n95), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[9]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n119) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n94), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[10]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n118) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n93), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[11]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n117) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n92), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[12]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n116) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n91), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[13]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n115) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_14_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n90), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[14]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n114) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_15_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n89), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[15]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n113) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_16_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n88), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[16]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n112) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_17_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n87), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[17]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n111) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_18_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n86), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_18_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n110) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_19_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n85), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_19_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n109) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_20_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n84), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_20_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n108) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_21_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n83), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_21_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n107) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_22_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n82), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_22_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n106) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_Q_int_reg_23_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n81), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_product_23_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_output_reg_n105) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U173 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n170), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n100) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U172 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n24), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n101) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U171 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n174), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n102) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U170 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n175), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n103) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U169 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n104) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U168 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n177), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n105) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U167 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n178), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n106) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U166 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n107) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U165 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n25), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n108) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U164 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n174), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n109) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U163 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n175), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n110) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U162 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n111) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U161 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n177), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n112) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U160 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n178), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n113) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U159 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n114) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U158 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op2_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n26), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n115) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U157 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n174), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n116) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U156 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n175), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n117) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U155 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n176), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n118) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U154 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n177), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n119) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U153 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n178), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n120) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U152 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n36), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n181) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U151 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n21), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n180) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U150 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n181), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n180), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n41) );
  XNOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U149 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n180), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n181), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n42) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U148 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op2_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op1_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n73) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U147 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n74) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U146 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n75) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U145 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n76) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U144 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n77) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U143 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n78) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U142 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n79) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U141 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n21), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n80) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U140 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n174), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n81) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U139 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n175), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n82) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U138 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n83) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U137 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n178), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n85) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U136 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n86) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U135 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n22), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n87) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U134 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n174), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n88) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U133 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n169), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n175), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n89) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U132 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n90) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U131 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n177), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n91) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U130 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n178), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n92) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U129 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n93) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U128 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_op2_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n94) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U127 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n174), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n95) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U126 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n176), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n97) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U125 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n177), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n98) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U124 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n178), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n99) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U123 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n179), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[0]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U122 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n21), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n168) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U121 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n175) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U120 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n177) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U119 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n170) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U118 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n25), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n172) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U117 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n24), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n171) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U116 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n22), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n169) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U115 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n174) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U114 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n176) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U113 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n178) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U112 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n179) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U111 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_n26), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n173) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U110 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[13]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U44 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n113), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n119), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n71), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n72) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U43 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n100), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n106), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n69), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n70) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U42 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n112), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n118), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n71), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n67), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n68) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U41 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n93), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n99), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n65), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n66) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U40 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n105), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n117), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n111), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n63), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n64) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U39 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n66), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n69), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n67), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n61), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n62) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U38 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n86), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n92), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n59), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n60) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U37 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n98), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n116), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n104), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n57), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n58) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U36 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n65), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n110), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n60), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n55), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n56) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U35 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n58), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n63), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n56), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n53), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n54) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U34 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n97), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n91), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n51), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n52) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U33 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n85), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n103), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n109), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n49), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n50) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U32 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n79), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n115), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n59), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n47), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n48) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U31 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n57), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n52), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n50), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n45), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n46) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U30 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n48), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n55), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n46), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n43), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n44) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U27 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n102), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n90), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n108), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n39), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n40) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n51), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n78), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n42), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n37), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n38) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U25 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n47), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n49), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n40), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n35), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n36) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U24 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n45), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n38), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n36), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n33), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n34) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U23 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n83), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n89), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n95), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n31), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n32) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U22 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n77), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n101), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n41), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n29), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n30) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U21 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n32), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n39), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n37), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n27), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n28) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U20 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n35), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n30), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n28), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n25), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n26) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U19 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n82), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n88), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n94), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n23), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n24) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U18 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n31), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n76), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n29), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n21), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n22) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U17 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n27), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n24), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n22), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n19), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n20) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U16 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n87), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n81), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n75), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n17), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n18) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U15 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n18), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n23), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n21), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n15), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n16) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U14 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n74), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n80), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n17), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n13), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n14) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n120), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n114), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n12), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[1]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U12 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n12), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n107), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n72), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n11), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[2]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n11), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n70), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n68), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n10), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[3]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n62), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n64), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n10), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n9), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[4]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n54), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n61), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n9), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n8), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[5]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n44), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n53), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n8), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n7), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[6]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n34), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n43), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n7), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n6), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[7]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U6 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n26), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n33), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n6), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n5), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[8]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n20), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n25), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n5), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n4), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[9]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n16), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n19), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n4), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n3), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[10]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n15), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n14), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n3), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n2), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[11]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_U2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n13), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n73), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n2), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_47_n1), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_2_mult_int[12]) );
  NOR3_X4 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U103 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_int_LE), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_), .A3(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n113), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U102 ( .A1(1'b0), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op2_int_6_) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U101 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_11_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_5_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n119) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U100 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n119), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n28) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U99 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_10_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_4_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n118) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U98 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n118), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n29) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U97 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_9_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_3_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n117) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U96 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n117), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n30) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U95 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_8_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_2_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n116) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U94 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n116), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n31) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U93 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_7_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_1_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n115) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U92 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n115), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n32) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U91 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_0_), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n114) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U90 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n114), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n33) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U89 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_11_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_5_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n126) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U88 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n126), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n10) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U87 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_10_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n124) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U86 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n124), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n12) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U85 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_9_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_3_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n123) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U84 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n123), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n14) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U83 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_8_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_2_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n122) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U82 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n122), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n16) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U81 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_7_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n121) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U80 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n121), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n18) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U79 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_6_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n120) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U78 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n120), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n20) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U77 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__1_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n153) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U76 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n153), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n39) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U75 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__0_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n152) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U74 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n152), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n40) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U73 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__3_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n155) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U72 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n155), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n37) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U71 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_25_), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n143), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_N35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n145) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U70 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n145), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n1) );
  AOI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U69 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n41), .B2(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__5_), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n157) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U68 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n157), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n35) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U67 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__4_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n156) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U66 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n156), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n36) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U65 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_coord_comp_2__2_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n41), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n154) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U64 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n154), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n38) );
  AOI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U63 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n27), .B2(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[41]), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op1_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n151) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U62 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n151), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n21) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U61 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[40]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[46]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n150) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U60 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n150), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n22) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U59 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[38]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[44]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n148) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U58 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n148), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n24) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U57 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[37]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[43]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n147) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U56 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n147), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n25) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U55 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[36]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[42]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n146) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U54 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n146), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n26) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U53 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[39]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n27), .B1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[45]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n149) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U52 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n149), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n23) );
  OR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U51 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_n36), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_rst_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n113) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U50 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_24_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n140) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U49 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n2), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n140), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n112) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U48 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_23_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n139) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U47 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n3), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n139), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n111) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U46 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_22_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n138) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U45 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n4), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n138), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n110) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U44 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_21_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n137) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U43 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n5), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n137), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n109) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U42 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_20_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n136) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U41 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n6), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n136), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n108) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U40 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_19_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n135) );
  OAI211_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U39 ( .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n7), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n141), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n135), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n107) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U38 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out_samp[47]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op1_int_6_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U37 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n41) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U36 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_12_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n127) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U35 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n19) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U34 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n19), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n8), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n127), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n100) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U33 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_13_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n128) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U32 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_1_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n17) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U31 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n17), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n7), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n128), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n101) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U30 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_14_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n129) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U29 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_2_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n15) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U28 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n15), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n6), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n129), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n102) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U27 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_15_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n130) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_3_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n13) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U25 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n13), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n5), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n130), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n103) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U24 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_16_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n131) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U23 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_4_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n11) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U22 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n11), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n4), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n131), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n104) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U21 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_17_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n132) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U20 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_5_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n9) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U19 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n9), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n3), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n132), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n105) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U18 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_18_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n133) );
  OAI221_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U17 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n8), .C1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n134), .C2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n2), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n133), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n106) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U16 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n27) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U15 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n143), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n134) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U14 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n113), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n125) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U12 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_12_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n2) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_7_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n7) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_8_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n6) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_9_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n5) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_10_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n4) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_11_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n3) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U6 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_N35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n141) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U5 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n113), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n144), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n143) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n134), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n34) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_U3 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n143), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n27), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n142) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n33), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_0_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n32), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_1_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n31), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_2_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n30), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_3_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n29), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_4_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n28), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_5_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n20), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_6_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n18), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_7_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n16), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_8_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n14), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_9_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n12), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_10_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n10), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_11_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_19_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n107), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_19_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_20_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n108), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_20_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_21_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n109), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_21_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_22_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n110), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_22_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_23_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n111), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_23_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_24_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n112), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_24_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_25_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n1), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_25_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_18_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n106), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_18_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_17_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n105), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_17_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_16_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n104), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_16_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_15_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n103), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_15_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_14_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n102), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_14_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n101), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_13_) );
  DFF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n100), .CK(clk), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_12_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n2) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_U5 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n9), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n8), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_rst_0_) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_U4 ( 
        .A1(MULT1_VALID), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n10) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_U6 ( 
        .A(MULT1_VALID), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n6) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_U3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n10), 
        .B(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n9), 
        .Z(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n7) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_count_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n7), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_1_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n9) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_count_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n6), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_count_int_0_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_ctrl_sign_gen_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n2) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[0]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[0]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[1]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[2]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[3]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[4]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[5]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[6]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[7]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[8]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[9]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[10]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[11]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[11]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[12]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[12]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_Q_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[13]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1_sampling_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[13]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_12_), 
        .B(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[0]), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_0_) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_12_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_n1) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1_1 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[1]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_13_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_n1), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[2]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_1_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1_2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[2]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_14_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[2]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[3]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_2_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1_3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[3]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_15_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[3]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[4]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_3_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1_4 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[4]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_16_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[4]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[5]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_4_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1_5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[5]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_17_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[5]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[6]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_5_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1_6 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[6]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_18_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[6]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[7]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_6_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1_7 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[7]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_19_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[7]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[8]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_7_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1_8 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[8]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_20_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[8]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[9]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_8_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1_9 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[9]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_21_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[9]), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[10]), .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_9_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1_10 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[10]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_22_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[10]), .CO(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[11]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_10_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1_11 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[11]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_23_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[11]), .CO(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[12]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_11_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1_12 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[12]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_24_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[12]), .CO(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[13]), 
        .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_12_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_U1_13 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add1[13]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_25_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_pp_sum_add_19_carry[13]), .S(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_N35) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_int_LE_FF_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_int_LE_FF_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_int_LE_FF_Q_int_reg ( 
        .D(MULT1_VALID), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_int_LE_FF_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_int_LE) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_RST_FFX_1_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_RST_FFX_1_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_RST_FFX_1_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_rst_0_), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_RST_FFX_1_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_rst_1_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_RST_FFX_2_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_RST_FFX_2_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_RST_FFX_2_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_rst_1_), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_RST_FFX_2_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_RST_FFX_2_Q) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_result_LE_FF_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_result_LE_FF_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_result_LE_FF_Q_int_reg ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_SUM_rst_0_), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_result_LE_FF_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_result_LE) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U57 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U56 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U55 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_5_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n147) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U54 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n123), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n147), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n99) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U53 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_4_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n148) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U52 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n124), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n148), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n100) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U51 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_3_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n149) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U50 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n125), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n149), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n101) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U49 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_2_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n150) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U48 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n126), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n150), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n102) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U47 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_1_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n151) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U46 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n127), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n151), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n103) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U45 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_5_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n135) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U44 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n111), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n135), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n87) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U43 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_result_LE), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n74) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U42 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_result_LE), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n72) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U41 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n134) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U40 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n110), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n134), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n86) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U39 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_4_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n136) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U38 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n112), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n136), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n88) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U37 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_3_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n137) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U36 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n113), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n137), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n89) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U35 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_2_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n138) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U34 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n114), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n138), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n90) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U33 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_1_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n139) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U32 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n115), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n139), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n91) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U31 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_0_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n140) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U30 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n116), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n140), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n92) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U29 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_11_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n141) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U28 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n117), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n141), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n93) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U27 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_10_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n142) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U26 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n118), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n142), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n94) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U25 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_9_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n143) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U24 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n119), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n143), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n95) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U23 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_8_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n144) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U22 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n120), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n144), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n96) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U21 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_7_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n145) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U20 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n121), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n145), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n97) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U19 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_6_), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n146) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U18 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n122), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n146), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n98) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U17 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_int_0_), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n152) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U16 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n128), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n152), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n104) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U15 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_11_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n129) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U14 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n105), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n129), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n81) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U13 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_10_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n130) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U12 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n106), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n130), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n82) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U11 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_9_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n131) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U10 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n107), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n131), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n83) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U9 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_8_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n132) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U8 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n108), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n132), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n84) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U7 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_add_out_7_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n133) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U6 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n109), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78), .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n133), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n85) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n74), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n78) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n74), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n77) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n72), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n76) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_U2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n72), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n75) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n104), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[0]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n128) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n103), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[1]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n127) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n102), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[2]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n126) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n101), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[3]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n125) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n100), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[4]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n124) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n99), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[5]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n123) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n98), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[6]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n122) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n97), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[7]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n121) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n96), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[8]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n120) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n95), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[9]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n119) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n94), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[10]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n118) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n93), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n79), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[11]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n117) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n92), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[12]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n116) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n91), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[13]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n115) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_14_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n90), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[14]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n114) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_15_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n89), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[15]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n113) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_16_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n88), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[16]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n112) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_17_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n87), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[17]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n111) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_18_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n86), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_18_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n110) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_19_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n85), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_19_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n109) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_20_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n84), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_20_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n108) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_21_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n83), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_21_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n107) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_22_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n82), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_22_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n106) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_Q_int_reg_23_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n81), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n80), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_product_23_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_output_reg_n105) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U173 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n170), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n100) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U172 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n24), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n101) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U171 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n174), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n102) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U170 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n175), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n103) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U169 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n104) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U168 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n177), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n105) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U167 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n178), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n106) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U166 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n171), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n107) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U165 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n25), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n108) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U164 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n174), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n109) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U163 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n175), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n110) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U162 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n111) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U161 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n177), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n112) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U160 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n178), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n113) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U159 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n172), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n114) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U158 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op2_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n26), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n115) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U157 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n174), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n116) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U156 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n175), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n117) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U155 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n176), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n118) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U154 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n177), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n119) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U153 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n178), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n120) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U152 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n36), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n181) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U151 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n21), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n180) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U150 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n181), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n180), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n41) );
  XNOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U149 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n180), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n181), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n42) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U148 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op2_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op1_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n73) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U147 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n74) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U146 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n75) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U145 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n76) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U144 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n77) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U143 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n78) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U142 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op1_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n79) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U141 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n21), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n80) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U140 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n174), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n81) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U139 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n175), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n82) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U138 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n83) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U137 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n178), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n85) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U136 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n168), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n86) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U135 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n22), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op2_int_6_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n87) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U134 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n174), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n88) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U133 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n169), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n175), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n89) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U132 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n176), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n90) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U131 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n177), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n91) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U130 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n178), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n92) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U129 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n179), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n169), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n93) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U128 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_op2_int_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n94) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U127 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n174), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n95) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U126 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n176), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n97) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U125 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n177), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n98) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U124 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n170), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n178), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n99) );
  NOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U123 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n173), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n179), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[0]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U122 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n21), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n168) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U121 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n175) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U120 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n177) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U119 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n170) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U118 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n25), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n172) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U117 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n24), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n171) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U116 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n22), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n169) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U115 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n174) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U114 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n176) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U113 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n178) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U112 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n40), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n179) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U111 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_n26), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n173) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U110 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[13]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U44 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n113), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n119), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n71), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n72) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U43 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n100), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n106), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n69), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n70) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U42 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n112), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n118), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n71), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n67), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n68) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U41 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n93), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n99), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n65), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n66) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U40 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n105), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n117), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n111), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n63), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n64) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U39 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n66), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n69), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n67), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n61), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n62) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U38 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n86), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n92), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n59), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n60) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U37 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n98), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n116), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n104), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n57), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n58) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U36 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n65), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n110), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n60), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n55), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n56) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U35 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n58), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n63), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n56), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n53), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n54) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U34 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n97), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n91), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n51), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n52) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U33 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n85), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n103), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n109), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n49), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n50) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U32 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n79), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n115), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n59), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n47), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n48) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U31 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n57), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n52), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n50), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n45), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n46) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U30 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n48), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n55), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n46), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n43), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n44) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U27 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n102), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n90), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n108), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n39), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n40) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n51), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n78), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n42), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n37), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n38) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U25 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n47), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n49), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n40), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n35), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n36) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U24 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n45), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n38), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n36), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n33), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n34) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U23 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n83), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n89), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n95), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n31), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n32) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U22 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n77), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n101), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n41), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n29), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n30) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U21 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n32), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n39), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n37), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n27), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n28) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U20 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n35), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n30), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n28), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n25), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n26) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U19 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n82), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n88), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n94), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n23), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n24) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U18 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n31), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n76), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n29), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n21), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n22) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U17 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n27), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n24), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n22), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n19), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n20) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U16 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n87), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n81), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n75), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n17), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n18) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U15 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n18), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n23), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n21), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n15), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n16) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U14 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n74), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n80), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n17), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n13), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n14) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n120), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n114), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n12), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[1]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U12 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n12), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n107), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n72), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n11), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[2]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n11), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n70), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n68), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n10), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[3]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n62), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n64), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n10), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n9), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[4]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n54), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n61), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n9), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n8), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[5]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n44), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n53), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n8), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n7), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[6]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n34), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n43), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n7), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n6), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[7]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U6 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n26), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n33), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n6), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n5), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[8]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n20), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n25), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n5), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n4), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[9]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n16), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n19), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n4), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n3), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[10]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n15), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n14), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n3), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n2), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[11]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_U2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n13), .B(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n73), .CI(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n2), .CO(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_47_n1), .S(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_X_3_mult_int[12]) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U26 ( 
        .A1(extimating_unit_MV0_out_int[10]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n11) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U25 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n22), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n11), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n34) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U24 ( 
        .A1(extimating_unit_MV0_out_int[9]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n10) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U23 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n21), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n10), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n32) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U22 ( 
        .A1(extimating_unit_MV0_out_int[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n9) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U21 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n20), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n35), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n9), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n31) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U20 ( 
        .A1(extimating_unit_MV0_out_int[7]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n8) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U19 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n19), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n35), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n8), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n30) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U18 ( 
        .A1(extimating_unit_MV0_out_int[6]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n7) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U17 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n18), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n35), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n7), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n29) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U16 ( 
        .A1(extimating_unit_MV0_out_int[5]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n6) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U15 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n17), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n35), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n6), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n28) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U14 ( 
        .A1(extimating_unit_MV0_out_int[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n5) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U13 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n16), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n35), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n5), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n27) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U12 ( 
        .A1(extimating_unit_MV0_out_int[3]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n4) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U11 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n15), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n35), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n4), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n26) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U10 ( 
        .A1(extimating_unit_MV0_out_int[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n3) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U9 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n14), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n35), .A(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n3), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n25) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U8 ( .A1(
        extimating_unit_MV0_out_int[1]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n2) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U7 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n13), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n35), .A(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n2), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n24) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U6 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n35), .A2(
        extimating_unit_MV0_out_int[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n1) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U5 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n12), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n35), .A(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n1), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n23) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U4 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n36) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U3 ( .A(
        ADD3_MVin_LE), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n33) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_U2 ( .A(
        ADD3_MVin_LE), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n35) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n32), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[9]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n21) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n34), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[10]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n22) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n24), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[1]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n13) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n25), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[2]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n14) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n26), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[3]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n15) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n27), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[4]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n16) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n28), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[5]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n17) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n29), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[6]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n18) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n30), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[7]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n19) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n31), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[8]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n20) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n23), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[0]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_0_n12) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U26 ( 
        .A1(extimating_unit_MV0_out_int[21]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n59) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U25 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n48), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n59), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n37) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U24 ( 
        .A1(extimating_unit_MV0_out_int[20]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n60) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U23 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n49), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n60), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n38) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U22 ( 
        .A1(extimating_unit_MV0_out_int[19]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n61) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U21 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n50), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n35), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n61), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n39) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U20 ( 
        .A1(extimating_unit_MV0_out_int[18]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n62) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U19 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n51), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n35), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n62), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n40) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U18 ( 
        .A1(extimating_unit_MV0_out_int[17]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n63) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U17 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n52), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n35), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n63), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n41) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U16 ( 
        .A1(extimating_unit_MV0_out_int[16]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n64) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U15 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n53), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n35), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n64), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n42) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U14 ( 
        .A1(extimating_unit_MV0_out_int[15]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n65) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U13 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n54), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n35), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n65), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n43) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U12 ( 
        .A1(extimating_unit_MV0_out_int[14]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n66) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U11 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n55), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n35), 
        .A(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n66), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n44) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U10 ( 
        .A1(extimating_unit_MV0_out_int[13]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n67) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U9 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n56), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n35), .A(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n67), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n45) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U8 ( .A1(
        extimating_unit_MV0_out_int[12]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n68) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U7 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n57), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n35), .A(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n68), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n46) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U6 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n35), .A2(
        extimating_unit_MV0_out_int[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n69) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U5 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n58), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n35), .A(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n69), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n47) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U4 ( .A(
        extimating_unit_RST1_int), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n36) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U3 ( .A(
        ADD3_MVin_LE), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n33) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_U2 ( .A(
        ADD3_MVin_LE), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n35) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n47), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[11]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n58) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n46), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[12]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n57) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n45), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[13]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n56) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n44), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[14]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n55) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n43), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[15]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n54) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n42), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[16]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n53) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n41), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[17]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n52) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n40), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[18]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n51) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n39), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[19]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n50) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n38), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[20]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n49) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n37), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n36), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[21]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_MV0_hv_in_ADD3_reg_1_n48) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U92 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n53) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U91 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[21]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n52), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[17]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n39) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U90 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n39), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n77) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U89 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[17]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[17]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n45), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n28) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U88 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n28), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n54) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U87 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[16]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[21]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n49), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n11) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U86 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[15]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[21]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n49), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n12) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U85 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[14]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[21]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n49), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n13) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U84 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[13]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[20]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n49), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n14) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U83 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[12]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[19]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n48), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n15) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U82 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[11]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[18]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n48), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n16) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U81 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[10]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[17]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n48), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n17) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U80 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[9]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[16]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n52), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n2) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U79 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[15]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n51), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n3) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U78 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[7]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[14]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n51), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n4) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U77 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[6]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[13]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n51), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n5) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U76 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[5]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[12]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n51), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n6) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U75 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n78), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n1) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U74 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n78), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n40) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U73 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[0]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n47), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n18) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U72 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n18), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n92) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U71 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n77), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n43), .B1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[18]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n38) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U70 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n38), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n75) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U69 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[16]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[16]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n48), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n29) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U68 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n11), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n74) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U67 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n29), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n55) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U66 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[15]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[15]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n45), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n30) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U65 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n12), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n73) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U64 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n30), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n56) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U63 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[14]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[14]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n44), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n31) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U62 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n13), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n72) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U61 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n31), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n57) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U60 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[13]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[13]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n44), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n32) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U59 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n14), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n79) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U58 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n32), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n58) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U57 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[12]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[12]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n44), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n33) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U56 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n15), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n80) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U55 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n33), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n59) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U54 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[11]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[11]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n44), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n34) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U53 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n16), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n81) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U52 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n34), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n60) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U51 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[10]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[10]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n43), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n35) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U50 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n17), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n82) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U49 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n35), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n61) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U48 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[9]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[9]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n47), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n19) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U47 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n2), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n83) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U46 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n19), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n62) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U45 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[8]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n47), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n20) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U44 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n3), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n84) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U43 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n20), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n63) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U42 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[7]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[7]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n47), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n21) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U41 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n4), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n85) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U40 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n21), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n64) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U39 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[6]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[6]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n46), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n22) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U38 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n5), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n86) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U37 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n22), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n65) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U36 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[5]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[5]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n46), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n23) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U35 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n6), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n87) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U34 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n23), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n66) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U33 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[4]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n46), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n24) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U32 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n7), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n88) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U31 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n24), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n67) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U30 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[3]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n50), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n8) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U29 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n25), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n68) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U28 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n8), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n89) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U27 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n50), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n9) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n26), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n69) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U25 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n9), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n90) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U24 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n77), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n43), .B1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[19]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n37) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U23 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n76) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U22 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[1]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n50), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n10) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U21 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[2]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n45), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n26) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U20 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[1]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[1]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n45), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n27) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U19 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[0]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[0]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n43), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n36) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U18 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n36), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n71) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U17 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[11]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n50), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n7) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U16 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_1[3]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_3[3]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n46), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n25) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U15 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n40), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n48) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U14 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n40), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n49) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n44) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U12 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n47) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n40), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n51) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n27), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n70) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n10), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n91) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n45) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n46) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U6 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n40), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n50) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n43) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n40), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n52) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n52), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n42) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count_reg ( .D(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n41), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n53), .Q(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n78) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .B(ADD3_VALID), 
        .Z(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n41) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n92), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n71), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_0_) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n92), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n71), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_n1)
         );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_1 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n70), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n91), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_n1), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[2]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_1_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n69), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n90), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[2]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[3]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_2_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n68), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n89), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[3]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[4]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_3_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_4 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n67), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n88), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[4]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[5]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_4_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n66), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n87), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[5]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[6]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_5_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_6 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n65), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n86), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[6]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[7]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_6_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_7 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n64), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n85), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[7]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[8]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_7_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_8 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n63), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n84), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[8]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[9]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_8_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_9 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n62), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n83), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[9]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[10]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_9_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_10 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n61), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n82), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[10]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[11]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_10_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_11 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n60), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n81), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[11]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[12]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_11_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_12 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n59), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n80), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[12]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[13]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_12_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_13 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n58), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n79), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[13]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[14]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_13_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_14 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n57), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n72), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[14]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[15]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_14_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_15 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n56), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n73), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[15]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[16]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_15_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_16 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n55), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n74), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[16]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[17]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_16_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_17 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n54), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n77), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[17]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[18]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_17_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_18 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n54), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n75), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[18]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[19]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_18_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_U1_19 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n54), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_n76), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_partial_adder_add_19_carry[19]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_19_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_19_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_19_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[19]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_18_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_18_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[18]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_17_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_17_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[17]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_16_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_16_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[16]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_15_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_15_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[15]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_14_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_14_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[14]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_13_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[13]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_12_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[12]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_11_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[11]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_10_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_9_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_8_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_7_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_6_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_5_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_4_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_3_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_2_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_1_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_0_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_samp[0]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U48 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U47 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n62) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U46 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_count), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n60) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U45 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_3_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n4) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U44 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n24), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n66), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n4), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n44)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U43 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_2_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n3) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U42 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n23), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n66), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n3), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n43)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U41 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_1_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n2) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U40 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n22), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n66), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n2), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n42)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U39 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n66), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n1) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U38 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n21), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n1), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n41)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U37 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_14_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n15) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U36 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n35), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n15), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n55)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U35 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_13_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n14) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U34 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n34), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n14), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n54)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U33 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_12_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n13) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U32 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n33), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n13), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n53)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U31 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_11_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n12) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U30 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n32), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n12), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n52)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U29 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_10_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n11) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U28 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n31), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n11), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n51)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U27 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_9_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n10) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U26 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n30), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n10), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n50)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U25 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_8_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n9) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U24 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n29), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n9), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n49)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U23 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_7_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n8) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U22 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n28), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n8), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n48)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U21 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n7) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U20 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n27), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n7), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n47)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U19 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_5_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n6) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U18 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n26), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n6), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n46)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U17 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_4_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n5) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U16 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n25), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n5), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n45)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U15 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_19_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n20) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U14 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n40), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n20), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n61)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U13 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_18_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n19) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U12 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n39), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n19), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n59)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U11 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_17_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n18) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U10 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n38), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n18), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n58)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U9 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_16_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n17) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U8 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n37), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n17), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n57)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U7 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_add_out_15_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n16) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U6 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n36), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n16), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n56)
         );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n62), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n66) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n62), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n65) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n60), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n64) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_U2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n60), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n63) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_15_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n56), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[15]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n36) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_14_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n55), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[14]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n35) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n54), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[13]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n34) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n53), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[12]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n33) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n52), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[11]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n32) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n51), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[10]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n31) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n50), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[9]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n30) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n49), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[8]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n29) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n48), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[7]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n28) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n47), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[6]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n27) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n46), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[5]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n26) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n45), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[4]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n25) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n44), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[3]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n24) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n43), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[2]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n23) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n42), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[1]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n22) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n41), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[0]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n21) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_16_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n57), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[16]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n37) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_17_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n58), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[17]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n38) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_18_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n59), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[18]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n39) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_Q_int_reg_19_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n61), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[19]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_1_output_register_n40) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U92 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n53) );
  OAI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U91 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[10]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n52), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[17]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n95) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U90 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n95), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n56) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U89 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[17]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[17]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n45), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n106) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U88 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n106), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n74) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U87 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[16]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[10]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n49), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n123) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U86 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[15]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[10]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n49), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n122) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U85 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[14]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[10]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n49), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n121) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U84 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[13]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[9]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n49), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n120) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U83 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[12]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[8]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n48), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n119) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U82 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[11]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[7]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n48), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n118) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U81 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[10]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[6]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n48), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n117) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U80 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[9]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[5]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n52), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n132) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U79 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[4]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n51), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n131) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U78 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[7]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[3]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n51), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n130) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U77 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[6]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[2]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n51), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n129) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U76 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[5]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[1]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n51), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n128) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U75 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n93), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n1) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U74 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n93), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n40) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U73 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[0]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n47), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n116) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U72 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n116), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n73) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U71 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n56), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n43), .B1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[18]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n96) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U70 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n96), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n55) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U69 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[16]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[16]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n48), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n105) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U68 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n123), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n57) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U67 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n105), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n75) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U66 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[15]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[15]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n45), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n104) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U65 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n122), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n58) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U64 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n104), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n76) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U63 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[14]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[14]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n44), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n103) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U62 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n121), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n59) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U61 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n103), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n77) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U60 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[13]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[13]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n44), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n102) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U59 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n120), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n60) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U58 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n102), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n79) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U57 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[12]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[12]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n44), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n101) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U56 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n119), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n61) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U55 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n101), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n80) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U54 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[11]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[11]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n44), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n100) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U53 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n118), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n62) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U52 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n100), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n81) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U51 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[10]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[10]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n43), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n99) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U50 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n117), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n63) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U49 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n99), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n82) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U48 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[9]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[9]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n47), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n115) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U47 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n132), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n64) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U46 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n115), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n83) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U45 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[8]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n47), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n114) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U44 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n131), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n65) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U43 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n114), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n84) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U42 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[7]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[7]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n47), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n113) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U41 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n130), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n66) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U40 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n113), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n85) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U39 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[6]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[6]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n46), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n112) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U38 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n129), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n67) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U37 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n112), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n86) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U36 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[5]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[5]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n46), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n111) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U35 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n128), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n68) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U34 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n111), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n87) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U33 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[4]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n46), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n110) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U32 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n127), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n69) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U31 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n110), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n88) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U30 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[3]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n50), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n126) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U29 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n109), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n89) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U28 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n126), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n70) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U27 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n50), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n125) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n108), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n90) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U25 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n125), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n71) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U24 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n56), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n43), .B1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[19]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n97) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U23 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n97), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n54) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U22 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[1]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(1'b0), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n50), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n124) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U21 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[2]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[2]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n45), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n108) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U20 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[1]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[1]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n45), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n107) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U19 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[0]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[0]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n43), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n98) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U18 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n98), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n92) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U17 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MV0_in_ADD3_ext[0]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n50), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n127) );
  AOI22_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U16 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_2[3]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42), .B1(
        extimating_unit_Pixel_Retrieval_Unit_MULT1_out_0[3]), .B2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n46), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n109) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U15 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n40), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n48) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U14 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n40), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n49) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U13 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n44) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U12 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n47) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U11 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n40), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n51) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n107), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n91) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n124), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n72) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n45) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n46) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U6 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n40), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n50) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n43) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n40), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n52) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n52), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n42) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .B(ADD3_VALID), 
        .Z(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n94) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count_reg ( .D(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n94), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n53), .Q(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n93) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n73), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n92), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_0_) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n73), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n92), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_n1)
         );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_1 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n91), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n72), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_n1), 
        .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[2]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_1_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n90), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n71), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[2]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[3]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_2_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n89), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n70), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[3]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[4]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_3_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_4 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n88), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n69), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[4]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[5]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_4_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n87), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n68), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[5]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[6]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_5_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_6 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n86), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n67), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[6]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[7]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_6_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_7 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n85), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n66), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[7]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[8]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_7_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_8 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n84), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n65), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[8]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[9]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_8_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_9 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n83), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n64), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[9]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[10]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_9_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_10 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n82), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n63), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[10]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[11]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_10_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_11 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n81), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n62), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[11]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[12]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_11_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_12 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n80), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n61), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[12]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[13]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_12_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_13 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n79), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n60), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[13]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[14]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_13_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_14 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n77), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n59), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[14]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[15]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_14_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_15 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n76), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n58), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[15]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[16]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_15_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_16 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n75), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n57), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[16]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[17]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_16_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_17 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n74), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n56), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[17]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[18]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_17_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_18 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n74), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n55), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[18]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[19]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_18_) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_U1_19 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n74), .B(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_n54), .CI(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_partial_adder_add_19_carry[19]), .S(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_19_) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_0_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[0]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_1_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_2_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_3_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_4_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_5_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_6_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_7_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_8_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_9_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_10_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_11_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[11]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_12_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[12]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_13_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[13]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_14_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_14_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[14]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_15_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_15_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[15]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_16_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_16_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[16]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_17_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_17_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[17]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_18_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_18_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[18]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_Q_int_reg_19_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_19_), .CK(clk), 
        .RN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_sampling_n1), 
        .Q(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_samp[19]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U48 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U47 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n62) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U46 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_count), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n60) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U45 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_3_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n124) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U44 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n104), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n66), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n124), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n84)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U43 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_2_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n125) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U42 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n105), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n66), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n125), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n85)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U41 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_1_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n126) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U40 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n106), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n66), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n126), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n86)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U39 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n66), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n127) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U38 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n107), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n127), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n87)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U37 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_14_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n113) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U36 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n93), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n113), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n73)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U35 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_13_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n114) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U34 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n94), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n114), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n74)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U33 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_12_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n115) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U32 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n95), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n115), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n75)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U31 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_11_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n116) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U30 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n96), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n116), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n76)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U29 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_10_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n117) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U28 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n97), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n117), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n77)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U27 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_9_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n118) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U26 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n98), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n118), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n78)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U25 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_8_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n119) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U24 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n99), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n119), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n79)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U23 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_7_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n120) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U22 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n100), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n120), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n80)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U21 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_6_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n121) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U20 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n101), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n121), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n81)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U19 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_5_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n122) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U18 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n102), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n122), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n82)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U17 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_4_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n123) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U16 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n103), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n123), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n83)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U15 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_19_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n108) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U14 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n88), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n108), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n68)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U13 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_18_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n109) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U12 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n89), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n109), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n69)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U11 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_17_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n110) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U10 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n90), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n110), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n70)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U9 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_16_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n111) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U8 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n91), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n111), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n71)
         );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U7 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_add_out_15_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n112) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U6 ( 
        .B1(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n92), 
        .B2(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64), 
        .A(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n112), 
        .ZN(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n72)
         );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n62), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n66) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n62), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n65) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n60), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n64) );
  BUF_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_U2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n60), .Z(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n63) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n87), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[0]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n107) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n86), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[1]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n106) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n85), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[2]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n105) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n84), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[3]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n104) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n83), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[4]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n103) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n82), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[5]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n102) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n81), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[6]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n101) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n80), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[7]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n100) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n79), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[8]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n99) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n78), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[9]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n98) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n77), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[10]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n97) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n76), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[11]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n96) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n75), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[12]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n95) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_13_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n74), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[13]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n94) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_14_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n73), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[14]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n93) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_15_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n72), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[15]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n92) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_16_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n71), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[16]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n91) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_17_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n70), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[17]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n90) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_18_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n69), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[18]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n89) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_Q_int_reg_19_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n68), 
        .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n67), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[19]), .QN(
        extimating_unit_Pixel_Retrieval_Unit_ADD3_0_output_register_n88) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U29 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[13]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n7), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[5]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U28 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[12]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n6), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[4]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U27 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[11]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n5), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[3]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[10]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n2), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[2]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U25 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[9]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[1]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U24 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_N2), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[8]), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[0]) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U23 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n12), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[18]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n25) );
  XNOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U22 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[19]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n25), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[11]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U21 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[18]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n12), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[10]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U20 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[17]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n11), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[9]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U19 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[16]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n10), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[8]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U18 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[15]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n9), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[7]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U17 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[14]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n8), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[6]) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U16 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n11), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[17]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n12) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U15 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n10), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[16]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n11) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U14 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n9), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[15]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n10) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U13 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n8), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[14]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n9) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U12 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n7), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[13]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n8) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U11 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n6), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[12]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n7) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U10 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n5), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n6) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U9 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n2), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[10]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n5) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U8 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[9]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n2) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U7 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_N2), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n1) );
  NOR4_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U6 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n4), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[0]), .A3(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[2]), .A4(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[1]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n3) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[7]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n26) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U4 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n3), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n26), .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[19]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_N0) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U3 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_N0), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[7]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_N2) );
  OR4_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_U2 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[3]), .A3(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[6]), .A4(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v[5]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_v_round_n4) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U29 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[13]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n7), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[5]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U28 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[12]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n6), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[4]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U27 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[11]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n5), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[3]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U26 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[10]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n2), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[2]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U25 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[9]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n1), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[1]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U24 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_N2), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[8]), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[0]) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U23 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n12), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[18]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n25) );
  XNOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U22 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[19]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n25), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[11]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U21 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[18]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n12), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[10]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U20 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[17]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n11), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[9]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U19 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[16]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n10), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[8]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U18 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[15]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n9), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[7]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U17 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[14]), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n8), .Z(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[6]) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U16 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n11), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[17]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n12) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U15 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n10), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[16]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n11) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U14 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n9), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[15]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n10) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U13 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n8), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[14]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n9) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U12 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n7), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[13]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n8) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U11 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n6), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[12]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n7) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U10 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n5), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[11]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n6) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U9 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n2), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[10]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n5) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U8 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n1), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[9]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n2) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U7 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[8]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_N2), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n1) );
  NOR4_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U6 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n27), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[0]), .A3(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[2]), .A4(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[1]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n28) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[7]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n26) );
  OAI21_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U4 ( .B1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n28), .B2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n26), .A(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[19]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_N0) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U3 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_N0), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[7]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_N2) );
  OR4_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_U2 ( .A1(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[4]), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[3]), .A3(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[6]), .A4(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h[5]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_ex_h_round_n27) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[0]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[0]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[1]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[2]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[3]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[4]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[5]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_Q_int_reg_6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[6]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_Q_int_reg_7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[7]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_Q_int_reg_8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[8]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_Q_int_reg_9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[9]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_Q_int_reg_10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[10]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_Q_int_reg_11_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_tmp[11]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[11]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_Q_int_reg_0_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[0]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[0]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_Q_int_reg_1_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[1]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_Q_int_reg_2_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[2]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_Q_int_reg_3_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[3]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_Q_int_reg_4_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[4]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_Q_int_reg_5_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[5]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_Q_int_reg_6_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[6]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_Q_int_reg_7_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[7]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_Q_int_reg_8_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[8]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_Q_int_reg_9_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[9]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_Q_int_reg_10_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[10]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_Q_int_reg_11_ ( .D(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_tmp[11]), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h_REG_n1), .Q(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[11]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_x_0_), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[0]), .Z(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[0]) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U1 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_x_0_), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_h[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_n1) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U1_1 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_h[1]), .B(
        extimating_unit_Pixel_Retrieval_Unit_x_1_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_n1), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[2]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[1]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U1_2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_h[2]), .B(
        extimating_unit_Pixel_Retrieval_Unit_x_2_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[2]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[3]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[2]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U1_3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_h[3]), .B(
        extimating_unit_Pixel_Retrieval_Unit_x_3_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[3]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[4]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[3]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U1_4 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_h[4]), .B(
        extimating_unit_Pixel_Retrieval_Unit_x_4_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[4]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[5]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[4]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U1_5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_h[5]), .B(
        extimating_unit_Pixel_Retrieval_Unit_x_5_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[5]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[6]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[5]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U1_6 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_h[6]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[6]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[7]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[6]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U1_7 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_h[7]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[7]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[8]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[7]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U1_8 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_h[8]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[8]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[9]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[8]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U1_9 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_h[9]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[9]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[10]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[9]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U1_10 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_h[10]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[10]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[11]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[10]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U1_11 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_h[11]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[11]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[12]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[11]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_U1_12 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_h[11]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_calculator_add_19_carry[12]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[12]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_y_counter_U5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_y_counter_n2) );
  NAND2_X1 extimating_unit_Pixel_Retrieval_Unit_y_counter_U4 ( .A1(incrY), 
        .A2(extimating_unit_Pixel_Retrieval_Unit_y_count_out_0_), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_y_counter_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_y_counter_count_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y_counter_n5), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_y_counter_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y_count_out_1_), .QN(
        extimating_unit_Pixel_Retrieval_Unit_y_counter_n3) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_y_counter_count_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y_counter_n7), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_y_counter_n2), .Q(
        extimating_unit_Pixel_Retrieval_Unit_y_count_out_0_) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_y_counter_U6 ( .A(incrY), .B(
        extimating_unit_Pixel_Retrieval_Unit_y_count_out_0_), .Z(
        extimating_unit_Pixel_Retrieval_Unit_y_counter_n7) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_y_counter_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_y_counter_n1), .B(
        extimating_unit_Pixel_Retrieval_Unit_y_counter_n3), .Z(
        extimating_unit_Pixel_Retrieval_Unit_y_counter_n5) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_n3), .B(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[0]), .Z(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[0]) );
  AND2_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U1 ( 
        .A1(extimating_unit_Pixel_Retrieval_Unit_n3), .A2(
        extimating_unit_Pixel_Retrieval_Unit_MVr_v[0]), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_n1) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U1_1 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_v[1]), .B(
        extimating_unit_Pixel_Retrieval_Unit_y_short_1_), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_n1), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[2]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[1]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U1_2 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_v[2]), .B(
        extimating_unit_Pixel_Retrieval_Unit_n6), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[2]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[3]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[2]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U1_3 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_v[3]), .B(
        extimating_unit_Pixel_Retrieval_Unit_n1), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[3]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[4]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[3]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U1_4 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_v[4]), .B(
        extimating_unit_Pixel_Retrieval_Unit_n7), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[4]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[5]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[4]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U1_5 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_v[5]), .B(
        extimating_unit_Pixel_Retrieval_Unit_n8), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[5]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[6]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[5]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U1_6 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_v[6]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[6]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[7]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[6]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U1_7 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_v[7]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[7]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[8]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[7]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U1_8 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_v[8]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[8]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[9]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[8]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U1_9 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_v[9]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[9]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[10]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[9]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U1_10 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_v[10]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[10]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[11]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[10]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U1_11 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_v[11]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[11]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[12]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[11]) );
  FA_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_U1_12 ( 
        .A(extimating_unit_Pixel_Retrieval_Unit_MVr_v[11]), .B(1'b0), .CI(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_calculator_add_19_carry[12]), .S(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[12]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x_0_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_n1), .Q(
        RADDR_CurCu_x[0]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x_1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_n1), .Q(
        RADDR_CurCu_x[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x_2_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_n1), .Q(
        RADDR_CurCu_x[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x_3_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_n1), .Q(
        RADDR_CurCu_x[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x_4_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_n1), .Q(
        RADDR_CurCu_x[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_x_5_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_x_sampling_n1), .Q(
        RADDR_CurCu_x[5]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_n3), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_n1), .Q(
        RADDR_CurCu_y[0]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_y_short_1_), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_n1), .Q(
        RADDR_CurCu_y[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_n6), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_n1), .Q(
        RADDR_CurCu_y[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_n1), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_n1), .Q(
        RADDR_CurCu_y[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_n7), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_n1), .Q(
        RADDR_CurCu_y[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_n8), .CK(clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_CurCu_y_sampling_n1), .Q(
        RADDR_CurCu_y[5]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[12]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1), .Q(
        RADDR_RefCu_x[12]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[11]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1), .Q(
        RADDR_RefCu_x[11]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[10]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1), .Q(
        RADDR_RefCu_x[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[9]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1), .Q(
        RADDR_RefCu_x[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[8]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1), .Q(
        RADDR_RefCu_x[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[7]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1), .Q(
        RADDR_RefCu_x[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[6]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1), .Q(
        RADDR_RefCu_x[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[5]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1), .Q(
        RADDR_RefCu_x[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[4]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1), .Q(
        RADDR_RefCu_x[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[3]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1), .Q(
        RADDR_RefCu_x[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[2]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1), .Q(
        RADDR_RefCu_x[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[1]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1), .Q(
        RADDR_RefCu_x[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_tmp[0]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_x_sampling_n1), .Q(
        RADDR_RefCu_x[0]) );
  INV_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_U3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n37), .ZN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_Q_int_reg_0_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[0]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1), .Q(
        RADDR_RefCu_y[0]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_Q_int_reg_1_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[1]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1), .Q(
        RADDR_RefCu_y[1]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_Q_int_reg_2_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[2]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1), .Q(
        RADDR_RefCu_y[2]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_Q_int_reg_3_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[3]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1), .Q(
        RADDR_RefCu_y[3]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_Q_int_reg_4_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[4]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1), .Q(
        RADDR_RefCu_y[4]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_Q_int_reg_5_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[5]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1), .Q(
        RADDR_RefCu_y[5]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_Q_int_reg_6_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[6]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1), .Q(
        RADDR_RefCu_y[6]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_Q_int_reg_7_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[7]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1), .Q(
        RADDR_RefCu_y[7]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_Q_int_reg_8_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[8]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1), .Q(
        RADDR_RefCu_y[8]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_Q_int_reg_9_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[9]), .CK(clk), .RN(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1), .Q(
        RADDR_RefCu_y[9]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_Q_int_reg_10_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[10]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1), .Q(
        RADDR_RefCu_y[10]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_Q_int_reg_11_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[11]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1), .Q(
        RADDR_RefCu_y[11]) );
  DFFR_X1 extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_Q_int_reg_12_ ( 
        .D(extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_tmp[12]), .CK(
        clk), .RN(
        extimating_unit_Pixel_Retrieval_Unit_RADDR_RefCu_y_sampling_n1), .Q(
        RADDR_RefCu_y[12]) );
  XOR2_X1 extimating_unit_Pixel_Retrieval_Unit_add_140_U1 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[11]), .B(
        extimating_unit_Pixel_Retrieval_Unit_n39), .Z(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[11]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_add_140_U1_1_1 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n59), .B(
        extimating_unit_Pixel_Retrieval_Unit_n60), .CO(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[2]), .S(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[1]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_add_140_U1_1_2 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n57), .B(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[2]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[3]), .S(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[2]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_add_140_U1_1_3 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n55), .B(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[3]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[4]), .S(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[3]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_add_140_U1_1_4 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n53), .B(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[4]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[5]), .S(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[4]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_add_140_U1_1_5 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n51), .B(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[5]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[6]), .S(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[5]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_add_140_U1_1_6 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n49), .B(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[6]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[7]), .S(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[6]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_add_140_U1_1_7 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n47), .B(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[7]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[8]), .S(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[7]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_add_140_U1_1_8 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n45), .B(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[8]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[9]), .S(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[8]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_add_140_U1_1_9 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n43), .B(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[9]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[10]), .S(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[9]) );
  HA_X1 extimating_unit_Pixel_Retrieval_Unit_add_140_U1_1_10 ( .A(
        extimating_unit_Pixel_Retrieval_Unit_n41), .B(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[10]), .CO(
        extimating_unit_Pixel_Retrieval_Unit_add_140_carry[11]), .S(
        extimating_unit_Pixel_Retrieval_Unit_R_SH2_out2_inv[10]) );
  INV_X1 extimating_unit_extimator_CU_U92 ( .A(RST), .ZN(
        extimating_unit_extimator_CU_n1) );
  INV_X1 extimating_unit_extimator_CU_U91 ( .A(
        extimating_unit_extimator_CU_last_block_x_int), .ZN(
        extimating_unit_extimator_CU_n3) );
  INV_X1 extimating_unit_extimator_CU_U90 ( .A(
        extimating_unit_extimator_CU_VALID_int), .ZN(
        extimating_unit_extimator_CU_n2) );
  AOI21_X1 extimating_unit_extimator_CU_U89 ( .B1(
        extimating_unit_extimator_CU_n23), .B2(eCU_PS[4]), .A(
        extimating_unit_extimator_CU_n38), .ZN(
        extimating_unit_extimator_CU_n37) );
  NAND4_X1 extimating_unit_extimator_CU_U88 ( .A1(
        extimating_unit_extimator_CU_n34), .A2(
        extimating_unit_extimator_CU_n35), .A3(
        extimating_unit_extimator_CU_n36), .A4(
        extimating_unit_extimator_CU_n37), .ZN(
        extimating_unit_SAD_tmp_RST_CU_int) );
  INV_X1 extimating_unit_extimator_CU_U87 ( .A(extimating_unit_CE_REPy_int), 
        .ZN(extimating_unit_extimator_CU_n5) );
  OAI21_X1 extimating_unit_extimator_CU_U86 ( .B1(eCU_PS[4]), .B2(
        extimating_unit_extimator_CU_n96), .A(extimating_unit_extimator_CU_n5), 
        .ZN(extimating_unit_CE_REPx_int) );
  INV_X1 extimating_unit_extimator_CU_U85 ( .A(
        extimating_unit_extimator_CU_n60), .ZN(extimating_unit_extimator_CU_n6) );
  AOI22_X1 extimating_unit_extimator_CU_U84 ( .A1(
        extimating_unit_extimator_CU_n56), .A2(
        extimating_unit_extimator_CU_n57), .B1(
        extimating_unit_extimator_CU_CountTerm_OUT_int), .B2(
        extimating_unit_extimator_CU_n15), .ZN(
        extimating_unit_extimator_CU_n50) );
  AND4_X1 extimating_unit_extimator_CU_U83 ( .A1(
        extimating_unit_extimator_CU_n52), .A2(
        extimating_unit_extimator_CU_n53), .A3(
        extimating_unit_extimator_CU_n54), .A4(
        extimating_unit_extimator_CU_n55), .ZN(
        extimating_unit_extimator_CU_n51) );
  NAND4_X1 extimating_unit_extimator_CU_U82 ( .A1(
        extimating_unit_extimator_CU_n6), .A2(extimating_unit_extimator_CU_n7), 
        .A3(extimating_unit_extimator_CU_n50), .A4(
        extimating_unit_extimator_CU_n51), .ZN(
        extimating_unit_extimator_CU_N182) );
  AOI21_X1 extimating_unit_extimator_CU_U81 ( .B1(
        extimating_unit_extimator_CU_n28), .B2(
        extimating_unit_extimator_CU_n57), .A(extimating_unit_extimator_CU_n23), .ZN(extimating_unit_extimator_CU_n82) );
  INV_X1 extimating_unit_extimator_CU_U80 ( .A(
        extimating_unit_extimator_CU_n82), .ZN(
        extimating_unit_extimator_CU_n13) );
  INV_X1 extimating_unit_extimator_CU_U79 ( .A(
        extimating_unit_extimator_CU_CountTerm_OUT_int), .ZN(
        extimating_unit_extimator_CU_n4) );
  NOR3_X1 extimating_unit_extimator_CU_U78 ( .A1(
        extimating_unit_extimator_CU_n73), .A2(
        extimating_unit_extimator_CU_n68), .A3(
        extimating_unit_extimator_CU_n74), .ZN(
        extimating_unit_extimator_CU_n72) );
  NOR3_X1 extimating_unit_extimator_CU_U77 ( .A1(
        extimating_unit_extimator_CU_n21), .A2(
        extimating_unit_extimator_CU_n67), .A3(OUT_LE), .ZN(
        extimating_unit_extimator_CU_n71) );
  NAND4_X1 extimating_unit_extimator_CU_U76 ( .A1(
        extimating_unit_extimator_CU_n70), .A2(
        extimating_unit_extimator_CU_n53), .A3(
        extimating_unit_extimator_CU_n71), .A4(
        extimating_unit_extimator_CU_n72), .ZN(
        extimating_unit_extimator_CU_N180) );
  NOR4_X1 extimating_unit_extimator_CU_U75 ( .A1(INTER_DATA_VALID_RESET), .A2(
        extimating_unit_extimator_CU_n49), .A3(
        extimating_unit_extimator_CU_n17), .A4(
        extimating_unit_extimator_CU_n22), .ZN(
        extimating_unit_extimator_CU_n64) );
  AOI21_X1 extimating_unit_extimator_CU_U74 ( .B1(
        extimating_unit_extimator_CU_last_cand_int), .B2(
        extimating_unit_extimator_CU_n67), .A(extimating_unit_extimator_CU_n68), .ZN(extimating_unit_extimator_CU_n63) );
  NAND4_X1 extimating_unit_extimator_CU_U73 ( .A1(
        extimating_unit_extimator_CU_n69), .A2(eCU_PS[1]), .A3(
        extimating_unit_extimator_CU_n28), .A4(
        extimating_unit_extimator_CU_n24), .ZN(
        extimating_unit_extimator_CU_n61) );
  NAND4_X1 extimating_unit_extimator_CU_U72 ( .A1(
        extimating_unit_extimator_CU_n61), .A2(
        extimating_unit_extimator_CU_n62), .A3(
        extimating_unit_extimator_CU_n63), .A4(
        extimating_unit_extimator_CU_n64), .ZN(
        extimating_unit_extimator_CU_N181) );
  AND3_X1 extimating_unit_extimator_CU_U71 ( .A1(
        extimating_unit_extimator_CU_last_block_x_int), .A2(
        extimating_unit_extimator_CU_n48), .A3(
        extimating_unit_extimator_CU_last_block_y_int), .ZN(
        extimating_unit_extimator_CU_n67) );
  NAND2_X1 extimating_unit_extimator_CU_U70 ( .A1(
        extimating_unit_extimator_CU_n89), .A2(eCU_PS[2]), .ZN(
        extimating_unit_extimator_CU_n96) );
  AND3_X1 extimating_unit_extimator_CU_U69 ( .A1(eCU_PS[2]), .A2(eCU_PS[1]), 
        .A3(extimating_unit_extimator_CU_n66), .ZN(
        extimating_unit_extimator_CU_n48) );
  NAND2_X1 extimating_unit_extimator_CU_U68 ( .A1(eCU_PS[3]), .A2(
        extimating_unit_extimator_CU_n24), .ZN(
        extimating_unit_extimator_CU_n41) );
  OAI21_X1 extimating_unit_extimator_CU_U67 ( .B1(
        extimating_unit_extimator_CU_Second_ready_int), .B2(
        extimating_unit_extimator_CU_n33), .A(extimating_unit_extimator_CU_n45), .ZN(extimating_unit_extimator_CU_n91) );
  AOI21_X1 extimating_unit_extimator_CU_U66 ( .B1(
        extimating_unit_extimator_CU_n15), .B2(extimating_unit_extimator_CU_n4), .A(extimating_unit_extimator_CU_n78), .ZN(extimating_unit_extimator_CU_n77)
         );
  NAND4_X1 extimating_unit_extimator_CU_U65 ( .A1(
        extimating_unit_extimator_CU_n75), .A2(
        extimating_unit_extimator_CU_n55), .A3(
        extimating_unit_extimator_CU_n76), .A4(
        extimating_unit_extimator_CU_n77), .ZN(
        extimating_unit_extimator_CU_n68) );
  NOR2_X1 extimating_unit_extimator_CU_U64 ( .A1(
        extimating_unit_extimator_CU_n28), .A2(
        extimating_unit_extimator_CU_n24), .ZN(
        extimating_unit_extimator_CU_n97) );
  NOR2_X1 extimating_unit_extimator_CU_U63 ( .A1(eCU_PS[1]), .A2(eCU_PS[0]), 
        .ZN(extimating_unit_extimator_CU_n89) );
  AOI22_X1 extimating_unit_extimator_CU_U62 ( .A1(
        extimating_unit_extimator_CU_n13), .A2(
        extimating_unit_extimator_CU_n25), .B1(eCU_PS[2]), .B2(
        extimating_unit_extimator_CU_n24), .ZN(
        extimating_unit_extimator_CU_n42) );
  NOR2_X1 extimating_unit_extimator_CU_U61 ( .A1(
        extimating_unit_extimator_CU_n41), .A2(
        extimating_unit_extimator_CU_n30), .ZN(
        extimating_unit_extimator_CU_n66) );
  NOR2_X1 extimating_unit_extimator_CU_U59 ( .A1(
        extimating_unit_extimator_CU_n30), .A2(eCU_PS[3]), .ZN(
        extimating_unit_extimator_CU_n69) );
  NAND4_X1 extimating_unit_extimator_CU_U58 ( .A1(
        extimating_unit_extimator_CU_n41), .A2(
        extimating_unit_extimator_CU_n36), .A3(
        extimating_unit_extimator_CU_n42), .A4(
        extimating_unit_extimator_CU_n43), .ZN(
        extimating_unit_RF_Addr_CU_int[0]) );
  NOR3_X1 extimating_unit_extimator_CU_U57 ( .A1(eCU_PS[3]), .A2(eCU_PS[4]), 
        .A3(extimating_unit_extimator_CU_n28), .ZN(
        extimating_unit_extimator_CU_n56) );
  AND2_X1 extimating_unit_extimator_CU_U56 ( .A1(
        extimating_unit_extimator_CU_n79), .A2(
        extimating_unit_extimator_CU_n30), .ZN(
        extimating_unit_extimator_CU_n90) );
  AND2_X1 extimating_unit_extimator_CU_U55 ( .A1(
        extimating_unit_extimator_CU_n92), .A2(
        extimating_unit_extimator_CU_n28), .ZN(
        extimating_unit_extimator_CU_n88) );
  NOR2_X1 extimating_unit_extimator_CU_U54 ( .A1(
        extimating_unit_extimator_CU_n29), .A2(eCU_PS[0]), .ZN(
        extimating_unit_extimator_CU_n92) );
  NOR2_X1 extimating_unit_extimator_CU_U53 ( .A1(
        extimating_unit_extimator_CU_n30), .A2(
        extimating_unit_extimator_CU_n29), .ZN(
        extimating_unit_extimator_CU_n57) );
  NOR2_X1 extimating_unit_extimator_CU_U52 ( .A1(eCU_PS[2]), .A2(eCU_PS[1]), 
        .ZN(extimating_unit_extimator_CU_n79) );
  NOR2_X1 extimating_unit_extimator_CU_U51 ( .A1(
        extimating_unit_extimator_CU_n24), .A2(
        extimating_unit_extimator_CU_n25), .ZN(
        extimating_unit_extimator_CU_n80) );
  OAI21_X1 extimating_unit_extimator_CU_U50 ( .B1(
        extimating_unit_extimator_CU_n57), .B2(eCU_PS[2]), .A(
        extimating_unit_extimator_CU_n80), .ZN(
        extimating_unit_extimator_CU_n98) );
  NAND2_X1 extimating_unit_extimator_CU_U49 ( .A1(
        extimating_unit_extimator_CU_n40), .A2(
        extimating_unit_extimator_CU_n39), .ZN(extimating_unit_RST_BLKx_int)
         );
  INV_X1 extimating_unit_extimator_CU_U48 ( .A(
        extimating_unit_extimator_CU_n39), .ZN(extimating_unit_RST_BLKy_int)
         );
  INV_X1 extimating_unit_extimator_CU_U47 ( .A(
        extimating_unit_extimator_CU_n33), .ZN(ADD3_MVin_LE_nSET) );
  NAND2_X1 extimating_unit_extimator_CU_U46 ( .A1(
        extimating_unit_extimator_CU_n81), .A2(
        extimating_unit_extimator_CU_n34), .ZN(CountTerm_EN) );
  INV_X1 extimating_unit_extimator_CU_U45 ( .A(extimating_unit_VALID_int), 
        .ZN(extimating_unit_extimator_CU_n31) );
  OAI22_X1 extimating_unit_extimator_CU_U44 ( .A1(
        extimating_unit_extimator_CU_n45), .A2(extimating_unit_extimator_CU_n2), .B1(extimating_unit_extimator_CU_n36), .B2(extimating_unit_extimator_CU_n31), 
        .ZN(extimating_unit_extimator_CU_n73) );
  INV_X1 extimating_unit_extimator_CU_U43 ( .A(
        extimating_unit_extimator_CU_n54), .ZN(
        extimating_unit_extimator_CU_n17) );
  NAND2_X1 extimating_unit_extimator_CU_U42 ( .A1(
        extimating_unit_extimator_CU_n27), .A2(
        extimating_unit_extimator_CU_n90), .ZN(
        extimating_unit_extimator_CU_n95) );
  NAND2_X1 extimating_unit_extimator_CU_U41 ( .A1(
        extimating_unit_extimator_CU_n90), .A2(
        extimating_unit_extimator_CU_n80), .ZN(
        extimating_unit_extimator_CU_n58) );
  NAND2_X1 extimating_unit_extimator_CU_U40 ( .A1(
        extimating_unit_extimator_CU_n27), .A2(
        extimating_unit_extimator_CU_n88), .ZN(
        extimating_unit_extimator_CU_n52) );
  AND2_X1 extimating_unit_extimator_CU_U39 ( .A1(
        extimating_unit_extimator_CU_n56), .A2(
        extimating_unit_extimator_CU_n92), .ZN(
        extimating_unit_extimator_CU_n78) );
  INV_X1 extimating_unit_extimator_CU_U38 ( .A(
        extimating_unit_extimator_CU_n81), .ZN(
        extimating_unit_extimator_CU_n21) );
  NOR3_X1 extimating_unit_extimator_CU_U37 ( .A1(
        extimating_unit_extimator_CU_n48), .A2(
        extimating_unit_extimator_CU_n49), .A3(
        extimating_unit_extimator_CU_n15), .ZN(
        extimating_unit_extimator_CU_n47) );
  NAND2_X1 extimating_unit_extimator_CU_U36 ( .A1(
        extimating_unit_extimator_CU_n66), .A2(
        extimating_unit_extimator_CU_n79), .ZN(
        extimating_unit_extimator_CU_n53) );
  NAND2_X1 extimating_unit_extimator_CU_U35 ( .A1(
        extimating_unit_extimator_CU_n88), .A2(
        extimating_unit_extimator_CU_n80), .ZN(
        extimating_unit_extimator_CU_n44) );
  INV_X1 extimating_unit_extimator_CU_U34 ( .A(
        extimating_unit_extimator_CU_n74), .ZN(
        extimating_unit_extimator_CU_n12) );
  AOI21_X1 extimating_unit_extimator_CU_U33 ( .B1(
        extimating_unit_extimator_CU_n15), .B2(extimating_unit_extimator_CU_n4), .A(extimating_unit_extimator_CU_n60), .ZN(extimating_unit_extimator_CU_n83)
         );
  AOI221_X1 extimating_unit_extimator_CU_U32 ( .B1(
        extimating_unit_extimator_CU_n48), .B2(extimating_unit_extimator_CU_n3), .C1(extimating_unit_extimator_CU_n91), .C2(extimating_unit_extimator_CU_n2), 
        .A(extimating_unit_extimator_CU_n78), .ZN(
        extimating_unit_extimator_CU_n84) );
  NAND4_X1 extimating_unit_extimator_CU_U31 ( .A1(
        extimating_unit_extimator_CU_n83), .A2(
        extimating_unit_extimator_CU_n12), .A3(
        extimating_unit_extimator_CU_n84), .A4(
        extimating_unit_extimator_CU_n85), .ZN(
        extimating_unit_extimator_CU_N179) );
  INV_X1 extimating_unit_extimator_CU_U30 ( .A(
        extimating_unit_extimator_CU_n96), .ZN(
        extimating_unit_extimator_CU_n23) );
  NAND2_X1 extimating_unit_extimator_CU_U29 ( .A1(
        extimating_unit_extimator_CU_n58), .A2(
        extimating_unit_extimator_CU_n59), .ZN(
        extimating_unit_extimator_CU_n38) );
  INV_X1 extimating_unit_extimator_CU_U28 ( .A(
        extimating_unit_extimator_CU_n41), .ZN(
        extimating_unit_extimator_CU_n27) );
  NAND2_X1 extimating_unit_extimator_CU_U27 ( .A1(
        extimating_unit_extimator_CU_n56), .A2(
        extimating_unit_extimator_CU_n89), .ZN(
        extimating_unit_extimator_CU_n62) );
  INV_X1 extimating_unit_extimator_CU_U26 ( .A(
        extimating_unit_extimator_CU_n59), .ZN(OUT_LE) );
  INV_X1 extimating_unit_extimator_CU_U25 ( .A(
        extimating_unit_extimator_CU_n94), .ZN(extimating_unit_CE_BLKx_int) );
  INV_X1 extimating_unit_extimator_CU_U24 ( .A(
        extimating_unit_extimator_CU_n45), .ZN(ADD3_MVin_LE_fSET) );
  INV_X1 extimating_unit_extimator_CU_U23 ( .A(
        extimating_unit_extimator_CU_n40), .ZN(extimating_unit_CE_BLKy_int) );
  OR2_X1 extimating_unit_extimator_CU_U22 ( .A1(ADD3_MVin_LE_fSET), .A2(
        extimating_unit_RST1_int), .ZN(extimating_unit_RST2_int) );
  NAND4_X1 extimating_unit_extimator_CU_U21 ( .A1(
        extimating_unit_extimator_CU_n52), .A2(
        extimating_unit_extimator_CU_n93), .A3(
        extimating_unit_extimator_CU_n40), .A4(
        extimating_unit_extimator_CU_n94), .ZN(
        extimating_unit_extimator_CU_n74) );
  INV_X1 extimating_unit_extimator_CU_U20 ( .A(
        extimating_unit_extimator_CU_n34), .ZN(
        extimating_unit_extimator_CU_n15) );
  NAND2_X1 extimating_unit_extimator_CU_U19 ( .A1(
        extimating_unit_extimator_CU_n33), .A2(
        extimating_unit_extimator_CU_n81), .ZN(INTER_DATA_VALID_RESET) );
  NOR2_X1 extimating_unit_extimator_CU_U18 ( .A1(
        extimating_unit_extimator_CU_n36), .A2(extimating_unit_VALID_int), 
        .ZN(extimating_unit_extimator_CU_n49) );
  INV_X1 extimating_unit_extimator_CU_U17 ( .A(
        extimating_unit_extimator_CU_n87), .ZN(extimating_unit_extimator_CU_n8) );
  NOR4_X1 extimating_unit_extimator_CU_U16 ( .A1(
        extimating_unit_extimator_CU_n86), .A2(eDONE), .A3(
        extimating_unit_extimator_CU_n8), .A4(extimating_unit_extimator_CU_n49), .ZN(extimating_unit_extimator_CU_n85) );
  OR2_X1 extimating_unit_extimator_CU_U15 ( .A1(INTER_DATA_VALID_SET), .A2(
        extimating_unit_RST1_int), .ZN(ADD3_MVin_LE_fRESET) );
  INV_X1 extimating_unit_extimator_CU_U14 ( .A(
        extimating_unit_extimator_CU_n93), .ZN(INTER_DATA_VALID_SET) );
  NOR2_X1 extimating_unit_extimator_CU_U13 ( .A1(eDONE), .A2(
        extimating_unit_RST2_int), .ZN(extimating_unit_extimator_CU_n35) );
  NOR2_X1 extimating_unit_extimator_CU_U12 ( .A1(INTER_DATA_VALID_RESET), .A2(
        extimating_unit_RST2_int), .ZN(extimating_unit_extimator_CU_n39) );
  NAND2_X1 extimating_unit_extimator_CU_U11 ( .A1(
        extimating_unit_extimator_CU_n27), .A2(
        extimating_unit_extimator_CU_n23), .ZN(
        extimating_unit_extimator_CU_n65) );
  INV_X1 extimating_unit_extimator_CU_U10 ( .A(
        extimating_unit_extimator_CU_n38), .ZN(extimating_unit_extimator_CU_n7) );
  NAND2_X1 extimating_unit_extimator_CU_U9 ( .A1(
        extimating_unit_extimator_CU_n7), .A2(extimating_unit_extimator_CU_n44), .ZN(extimating_unit_RF_Addr_CU_int[1]) );
  INV_X1 extimating_unit_extimator_CU_U8 ( .A(extimating_unit_extimator_CU_n44), .ZN(eDONE) );
  NAND2_X1 extimating_unit_extimator_CU_U7 ( .A1(
        extimating_unit_extimator_CU_n46), .A2(
        extimating_unit_extimator_CU_n95), .ZN(extimating_unit_CE_REPy_int) );
  NOR3_X1 extimating_unit_extimator_CU_U6 ( .A1(extimating_unit_CE_BLKx_int), 
        .A2(INTER_DATA_VALID_RESET), .A3(extimating_unit_CE_BLKy_int), .ZN(
        extimating_unit_extimator_CU_n46) );
  NOR4_X1 extimating_unit_extimator_CU_U5 ( .A1(
        extimating_unit_RF_Addr_CU_int[1]), .A2(extimating_unit_CE_REPy_int), 
        .A3(INTER_DATA_VALID_SET), .A4(extimating_unit_extimator_CU_n15), .ZN(
        extimating_unit_extimator_CU_n43) );
  INV_X1 extimating_unit_extimator_CU_U4 ( .A(extimating_unit_extimator_CU_n35), .ZN(extimating_unit_READY_RST_int) );
  INV_X1 extimating_unit_extimator_CU_U3 ( .A(extimating_unit_extimator_CU_n65), .ZN(extimating_unit_extimator_CU_n22) );
  DFFR_X1 extimating_unit_extimator_CU_PS_reg_1_ ( .D(eCU_NS[1]), .CK(clk), 
        .RN(extimating_unit_extimator_CU_n1), .Q(eCU_PS[1]), .QN(
        extimating_unit_extimator_CU_n29) );
  DFFR_X1 extimating_unit_extimator_CU_PS_reg_0_ ( .D(eCU_NS[0]), .CK(clk), 
        .RN(extimating_unit_extimator_CU_n1), .Q(eCU_PS[0]), .QN(
        extimating_unit_extimator_CU_n30) );
  DFFR_X1 extimating_unit_extimator_CU_PS_reg_2_ ( .D(eCU_NS[2]), .CK(clk), 
        .RN(extimating_unit_extimator_CU_n1), .Q(eCU_PS[2]), .QN(
        extimating_unit_extimator_CU_n28) );
  DFFR_X1 extimating_unit_extimator_CU_PS_reg_4_ ( .D(eCU_NS[4]), .CK(clk), 
        .RN(extimating_unit_extimator_CU_n1), .Q(eCU_PS[4]), .QN(
        extimating_unit_extimator_CU_n24) );
  DFFR_X1 extimating_unit_extimator_CU_PS_reg_3_ ( .D(eCU_NS[3]), .CK(clk), 
        .RN(extimating_unit_extimator_CU_n1), .Q(eCU_PS[3]), .QN(
        extimating_unit_extimator_CU_n25) );
  NAND3_X1 extimating_unit_extimator_CU_U112 ( .A1(
        extimating_unit_extimator_CU_n25), .A2(
        extimating_unit_extimator_CU_n24), .A3(
        extimating_unit_extimator_CU_n88), .ZN(
        extimating_unit_extimator_CU_n93) );
  NAND3_X1 extimating_unit_extimator_CU_U111 ( .A1(
        extimating_unit_extimator_CU_n25), .A2(
        extimating_unit_extimator_CU_n24), .A3(
        extimating_unit_extimator_CU_n90), .ZN(
        extimating_unit_extimator_CU_n87) );
  NAND3_X1 extimating_unit_extimator_CU_U110 ( .A1(
        extimating_unit_extimator_CU_n79), .A2(eCU_PS[4]), .A3(
        extimating_unit_extimator_CU_n69), .ZN(
        extimating_unit_extimator_CU_n94) );
  NAND3_X1 extimating_unit_extimator_CU_U109 ( .A1(eCU_PS[4]), .A2(
        extimating_unit_extimator_CU_n25), .A3(
        extimating_unit_extimator_CU_n88), .ZN(
        extimating_unit_extimator_CU_n33) );
  NAND3_X1 extimating_unit_extimator_CU_U108 ( .A1(
        extimating_unit_extimator_CU_n92), .A2(
        extimating_unit_extimator_CU_n25), .A3(
        extimating_unit_extimator_CU_n97), .ZN(
        extimating_unit_extimator_CU_n81) );
  NAND3_X1 extimating_unit_extimator_CU_U107 ( .A1(eCU_PS[4]), .A2(
        extimating_unit_extimator_CU_n25), .A3(
        extimating_unit_extimator_CU_n90), .ZN(
        extimating_unit_extimator_CU_n40) );
  NAND3_X1 extimating_unit_extimator_CU_U106 ( .A1(
        extimating_unit_extimator_CU_n69), .A2(eCU_PS[1]), .A3(
        extimating_unit_extimator_CU_n97), .ZN(
        extimating_unit_extimator_CU_n34) );
  NAND3_X1 extimating_unit_extimator_CU_U105 ( .A1(
        extimating_unit_extimator_CU_n79), .A2(
        extimating_unit_extimator_CU_n24), .A3(
        extimating_unit_extimator_CU_n69), .ZN(
        extimating_unit_extimator_CU_n45) );
  NAND3_X1 extimating_unit_extimator_CU_U104 ( .A1(
        extimating_unit_extimator_CU_n69), .A2(
        extimating_unit_extimator_CU_n29), .A3(
        extimating_unit_extimator_CU_n97), .ZN(
        extimating_unit_extimator_CU_n36) );
  NAND3_X1 extimating_unit_extimator_CU_U103 ( .A1(
        extimating_unit_extimator_CU_n45), .A2(
        extimating_unit_extimator_CU_n33), .A3(
        extimating_unit_extimator_CU_n36), .ZN(extimating_unit_LE_ab_CU_int)
         );
  NAND3_X1 extimating_unit_extimator_CU_U101 ( .A1(eCU_PS[2]), .A2(
        extimating_unit_extimator_CU_n92), .A3(
        extimating_unit_extimator_CU_n27), .ZN(
        extimating_unit_extimator_CU_n75) );
  NAND3_X1 extimating_unit_extimator_CU_U100 ( .A1(
        extimating_unit_extimator_CU_n65), .A2(
        extimating_unit_extimator_CU_n95), .A3(
        extimating_unit_extimator_CU_n75), .ZN(
        extimating_unit_extimator_CU_n60) );
  NAND3_X1 extimating_unit_extimator_CU_U99 ( .A1(
        extimating_unit_extimator_CU_n81), .A2(
        extimating_unit_extimator_CU_n58), .A3(
        extimating_unit_extimator_CU_n62), .ZN(
        extimating_unit_extimator_CU_n86) );
  NAND3_X1 extimating_unit_extimator_CU_U98 ( .A1(
        extimating_unit_extimator_CU_n13), .A2(
        extimating_unit_extimator_CU_n25), .A3(eCU_PS[4]), .ZN(
        extimating_unit_extimator_CU_n70) );
  NAND3_X1 extimating_unit_extimator_CU_U97 ( .A1(
        extimating_unit_extimator_CU_n79), .A2(
        extimating_unit_extimator_CU_n80), .A3(eCU_PS[0]), .ZN(
        extimating_unit_extimator_CU_n59) );
  NAND3_X1 extimating_unit_extimator_CU_U96 ( .A1(eCU_PS[2]), .A2(
        extimating_unit_extimator_CU_n29), .A3(
        extimating_unit_extimator_CU_n66), .ZN(
        extimating_unit_extimator_CU_n55) );
  NAND3_X1 extimating_unit_extimator_CU_U95 ( .A1(eCU_PS[0]), .A2(
        extimating_unit_extimator_CU_n29), .A3(
        extimating_unit_extimator_CU_n56), .ZN(
        extimating_unit_extimator_CU_n76) );
  NAND3_X1 extimating_unit_extimator_CU_U94 ( .A1(eCU_PS[1]), .A2(
        extimating_unit_extimator_CU_n28), .A3(
        extimating_unit_extimator_CU_n66), .ZN(
        extimating_unit_extimator_CU_n54) );
  NAND3_X1 extimating_unit_extimator_CU_U93 ( .A1(
        extimating_unit_extimator_CU_n46), .A2(extimating_unit_extimator_CU_n7), .A3(extimating_unit_extimator_CU_n47), .ZN(extimating_unit_extimator_CU_N183) );
  NAND2_X2 extimating_unit_extimator_CU_U60 ( .A1(
        extimating_unit_extimator_CU_n87), .A2(
        extimating_unit_extimator_CU_n98), .ZN(extimating_unit_RST1_int) );
  DLH_X1 extimating_unit_extimator_CU_NS_reg_4_ ( .G(1'b1), .D(
        extimating_unit_extimator_CU_N183), .Q(eCU_NS[4]) );
  DLH_X1 extimating_unit_extimator_CU_NS_reg_2_ ( .G(1'b1), .D(
        extimating_unit_extimator_CU_N181), .Q(eCU_NS[2]) );
  DLH_X1 extimating_unit_extimator_CU_NS_reg_3_ ( .G(1'b1), .D(
        extimating_unit_extimator_CU_N182), .Q(eCU_NS[3]) );
  DLH_X1 extimating_unit_extimator_CU_NS_reg_1_ ( .G(1'b1), .D(
        extimating_unit_extimator_CU_N180), .Q(eCU_NS[1]) );
  DLH_X1 extimating_unit_extimator_CU_NS_reg_0_ ( .G(1'b1), .D(
        extimating_unit_extimator_CU_N179), .Q(eCU_NS[0]) );
  INV_X1 extimating_unit_extimator_CU_VALID_samp_U3 ( .A(RST), .ZN(
        extimating_unit_extimator_CU_VALID_samp_n1) );
  DFFR_X1 extimating_unit_extimator_CU_VALID_samp_Q_int_reg ( .D(
        extimating_unit_VALID_int), .CK(clk), .RN(
        extimating_unit_extimator_CU_VALID_samp_n1), .Q(
        extimating_unit_extimator_CU_VALID_int) );
  INV_X1 extimating_unit_extimator_CU_last_block_x_samp_U3 ( .A(RST), .ZN(
        extimating_unit_extimator_CU_last_block_x_samp_n1) );
  DFFR_X1 extimating_unit_extimator_CU_last_block_x_samp_Q_int_reg ( .D(
        last_block_x), .CK(clk), .RN(
        extimating_unit_extimator_CU_last_block_x_samp_n1), .Q(
        extimating_unit_extimator_CU_last_block_x_int) );
  INV_X1 extimating_unit_extimator_CU_last_block_y_samp_U3 ( .A(RST), .ZN(
        extimating_unit_extimator_CU_last_block_y_samp_n1) );
  DFFR_X1 extimating_unit_extimator_CU_last_block_y_samp_Q_int_reg ( .D(
        last_block_y), .CK(clk), .RN(
        extimating_unit_extimator_CU_last_block_y_samp_n1), .Q(
        extimating_unit_extimator_CU_last_block_y_int) );
  INV_X1 extimating_unit_extimator_CU_last_cand_samp_U3 ( .A(RST), .ZN(
        extimating_unit_extimator_CU_last_cand_samp_n1) );
  DFFR_X1 extimating_unit_extimator_CU_last_cand_samp_Q_int_reg ( .D(last_cand), .CK(clk), .RN(extimating_unit_extimator_CU_last_cand_samp_n1), .Q(
        extimating_unit_extimator_CU_last_cand_int) );
  INV_X1 extimating_unit_extimator_CU_Second_ready_samp_U3 ( .A(RST), .ZN(
        extimating_unit_extimator_CU_Second_ready_samp_n1) );
  DFFR_X1 extimating_unit_extimator_CU_Second_ready_samp_Q_int_reg ( .D(
        Second_ready), .CK(clk), .RN(
        extimating_unit_extimator_CU_Second_ready_samp_n1), .Q(
        extimating_unit_extimator_CU_Second_ready_int) );
  INV_X1 extimating_unit_extimator_CU_CountTerm_OUT_samp_U3 ( .A(RST), .ZN(
        extimating_unit_extimator_CU_CountTerm_OUT_samp_n1) );
  DFFR_X1 extimating_unit_extimator_CU_CountTerm_OUT_samp_Q_int_reg ( .D(
        CountTerm_OUT), .CK(clk), .RN(
        extimating_unit_extimator_CU_CountTerm_OUT_samp_n1), .Q(
        extimating_unit_extimator_CU_CountTerm_OUT_int) );
  INV_X1 extimating_unit_Ready_Handler_U12 ( .A(RST), .ZN(
        extimating_unit_Ready_Handler_n1) );
  XNOR2_X1 extimating_unit_Ready_Handler_U11 ( .A(
        extimating_unit_Ready_Handler_n9), .B(
        extimating_unit_Ready_Handler_PS_1_), .ZN(
        extimating_unit_Ready_Handler_n8) );
  NOR2_X1 extimating_unit_Ready_Handler_U10 ( .A1(
        extimating_unit_Ready_Handler_PS_2_), .A2(
        extimating_unit_Ready_Handler_n8), .ZN(
        extimating_unit_Ready_Handler_NS[1]) );
  AND2_X1 extimating_unit_Ready_Handler_U9 ( .A1(
        extimating_unit_Ready_Handler_PS_0_), .A2(
        extimating_unit_Ready_Handler_n5), .ZN(eREADY) );
  AND2_X1 extimating_unit_Ready_Handler_U8 ( .A1(extimating_unit_VALID_int), 
        .A2(extimating_unit_Ready_Handler_PS_0_), .ZN(
        extimating_unit_Ready_Handler_n9) );
  AND2_X1 extimating_unit_Ready_Handler_U7 ( .A1(extimating_unit_READY_RST_int), .A2(extimating_unit_Ready_Handler_PS_0_), .ZN(
        extimating_unit_Ready_Handler_n6) );
  INV_X1 extimating_unit_Ready_Handler_U6 ( .A(Second_ready), .ZN(
        extimating_unit_Ready_Handler_n4) );
  OAI21_X1 extimating_unit_Ready_Handler_U5 ( .B1(
        extimating_unit_Ready_Handler_n6), .B2(
        extimating_unit_Ready_Handler_n4), .A(extimating_unit_Ready_Handler_n7), .ZN(extimating_unit_Ready_Handler_NS[2]) );
  NOR2_X1 extimating_unit_Ready_Handler_U4 ( .A1(
        extimating_unit_Ready_Handler_n5), .A2(
        extimating_unit_Ready_Handler_PS_1_), .ZN(Second_ready) );
  INV_X1 extimating_unit_Ready_Handler_U3 ( .A(
        extimating_unit_Ready_Handler_n9), .ZN(
        extimating_unit_Ready_Handler_n2) );
  DFFR_X1 extimating_unit_Ready_Handler_PS_reg_1_ ( .D(
        extimating_unit_Ready_Handler_NS[1]), .CK(clk), .RN(
        extimating_unit_Ready_Handler_n1), .Q(
        extimating_unit_Ready_Handler_PS_1_), .QN(
        extimating_unit_Ready_Handler_n3) );
  DFFR_X1 extimating_unit_Ready_Handler_PS_reg_2_ ( .D(
        extimating_unit_Ready_Handler_NS[2]), .CK(clk), .RN(
        extimating_unit_Ready_Handler_n1), .Q(
        extimating_unit_Ready_Handler_PS_2_), .QN(
        extimating_unit_Ready_Handler_n5) );
  NAND3_X1 extimating_unit_Ready_Handler_U13 ( .A1(
        extimating_unit_Ready_Handler_PS_1_), .A2(eREADY), .A3(
        extimating_unit_VALID_int), .ZN(extimating_unit_Ready_Handler_n7) );
  SDFFR_X1 extimating_unit_Ready_Handler_PS_reg_0_ ( .D(
        extimating_unit_Ready_Handler_n2), .SI(
        extimating_unit_Ready_Handler_n3), .SE(
        extimating_unit_Ready_Handler_PS_2_), .CK(clk), .RN(
        extimating_unit_Ready_Handler_n1), .Q(
        extimating_unit_Ready_Handler_PS_0_) );
  CLKBUF_X1 extimating_unit_CU_adapter_U19 ( .A(RST), .Z(
        extimating_unit_CU_adapter_n9) );
  INV_X1 extimating_unit_CU_adapter_U18 ( .A(clk), .ZN(
        extimating_unit_CU_adapter_n1) );
  BUF_X1 extimating_unit_CU_adapter_U17 ( .A(RST), .Z(
        extimating_unit_CU_adapter_n6) );
  BUF_X1 extimating_unit_CU_adapter_U16 ( .A(RST), .Z(
        extimating_unit_CU_adapter_n5) );
  BUF_X1 extimating_unit_CU_adapter_U15 ( .A(RST), .Z(
        extimating_unit_CU_adapter_n4) );
  BUF_X1 extimating_unit_CU_adapter_U14 ( .A(RST), .Z(
        extimating_unit_CU_adapter_n3) );
  BUF_X1 extimating_unit_CU_adapter_U13 ( .A(RST), .Z(
        extimating_unit_CU_adapter_n2) );
  INV_X1 extimating_unit_CU_adapter_U12 ( .A(INTER_DATA_VALID_SET), .ZN(
        extimating_unit_CU_adapter_n14) );
  INV_X1 extimating_unit_CU_adapter_U11 ( .A(
        extimating_unit_CU_adapter_MULT1_VALID_int_0_), .ZN(
        extimating_unit_CU_adapter_n10) );
  OAI21_X1 extimating_unit_CU_adapter_U10 ( .B1(
        extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_int[2]), .B2(
        extimating_unit_CU_adapter_n10), .A(extimating_unit_CU_adapter_n14), 
        .ZN(extimating_unit_CU_adapter_idv_sel) );
  INV_X1 extimating_unit_CU_adapter_U9 ( .A(ADD3_MVin_LE_fRESET), .ZN(
        extimating_unit_CU_adapter_n13) );
  NAND2_X1 extimating_unit_CU_adapter_U8 ( .A1(ADD3_MVin_LE_fSET), .A2(
        extimating_unit_CU_adapter_n13), .ZN(extimating_unit_CU_adapter_n8) );
  AOI21_X1 extimating_unit_CU_adapter_U7 ( .B1(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[9]), .B2(
        extimating_unit_CU_adapter_n13), .A(
        extimating_unit_CU_adapter_A3MVin_LE_samp), .ZN(
        extimating_unit_CU_adapter_n7) );
  NAND2_X1 extimating_unit_CU_adapter_U6 ( .A1(extimating_unit_CU_adapter_n7), 
        .A2(extimating_unit_CU_adapter_n8), .ZN(ADD3_MVin_LE) );
  INV_X1 extimating_unit_CU_adapter_U5 ( .A(extimating_unit_RF_Addr_CU_int[0]), 
        .ZN(extimating_unit_CU_adapter_n12) );
  INV_X1 extimating_unit_CU_adapter_U4 ( .A(BestCand), .ZN(
        extimating_unit_CU_adapter_n11) );
  AOI21_X1 extimating_unit_CU_adapter_U3 ( .B1(
        extimating_unit_RF_Addr_CU_int[1]), .B2(extimating_unit_CU_adapter_n11), .A(extimating_unit_CU_adapter_n12), .ZN(extimating_unit_RF_Addr_DP_int) );
  DFF_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_fRESET_half_delayed_reg ( .D(
        ADD3_MVin_LE_fRESET), .CK(extimating_unit_CU_adapter_n1), .Q(
        extimating_unit_CU_adapter_ADD3_MVin_LE_fRESET_half_delayed) );
  INV_X1 extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_delay_1_U3 ( .A(
        extimating_unit_CU_adapter_n2), .ZN(
        extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_delay_1_n1) );
  DFFR_X1 extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_delay_1_Q_int_reg ( 
        .D(INTER_DATA_VALID_RESET), .CK(clk), .RN(
        extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_delay_1_n1), .Q(
        extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_int[1]) );
  INV_X1 extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_delay_2_U3 ( .A(
        extimating_unit_CU_adapter_n2), .ZN(
        extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_delay_2_n1) );
  DFFR_X1 extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_delay_2_Q_int_reg ( 
        .D(extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_int[1]), .CK(clk), 
        .RN(extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_delay_2_n1), .Q(
        extimating_unit_CU_adapter_INTER_DATA_VALID_RESET_int[2]) );
  INV_X1 extimating_unit_CU_adapter_inter_data_valid_FlFl_U3 ( .A(
        extimating_unit_CU_adapter_n2), .ZN(
        extimating_unit_CU_adapter_inter_data_valid_FlFl_n1) );
  DFFR_X1 extimating_unit_CU_adapter_inter_data_valid_FlFl_Q_int_reg ( .D(
        extimating_unit_CU_adapter_idv_sel), .CK(clk), .RN(
        extimating_unit_CU_adapter_inter_data_valid_FlFl_n1), .Q(
        extimating_unit_CU_adapter_MULT1_VALID_int_0_) );
  INV_X1 extimating_unit_CU_adapter_MULT1_VALID_delay_1_U3 ( .A(
        extimating_unit_CU_adapter_n2), .ZN(
        extimating_unit_CU_adapter_MULT1_VALID_delay_1_n1) );
  DFFR_X1 extimating_unit_CU_adapter_MULT1_VALID_delay_1_Q_int_reg ( .D(
        extimating_unit_CU_adapter_MULT1_VALID_int_0_), .CK(clk), .RN(
        extimating_unit_CU_adapter_MULT1_VALID_delay_1_n1), .Q(
        extimating_unit_CU_adapter_MULT1_VALID_int_1_) );
  INV_X1 extimating_unit_CU_adapter_MULT1_VALID_delay_2_U3 ( .A(
        extimating_unit_CU_adapter_n2), .ZN(
        extimating_unit_CU_adapter_MULT1_VALID_delay_2_n1) );
  DFFR_X1 extimating_unit_CU_adapter_MULT1_VALID_delay_2_Q_int_reg ( .D(
        extimating_unit_CU_adapter_MULT1_VALID_int_1_), .CK(clk), .RN(
        extimating_unit_CU_adapter_MULT1_VALID_delay_2_n1), .Q(MULT1_VALID) );
  INV_X1 extimating_unit_CU_adapter_ADD3_VALID_delay_1_U3 ( .A(
        extimating_unit_CU_adapter_n2), .ZN(
        extimating_unit_CU_adapter_ADD3_VALID_delay_1_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_VALID_delay_1_Q_int_reg ( .D(
        MULT1_VALID), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_VALID_delay_1_n1), .Q(
        extimating_unit_CU_adapter_ADD3_VALID_int[1]) );
  INV_X1 extimating_unit_CU_adapter_ADD3_VALID_delay_2_U3 ( .A(
        extimating_unit_CU_adapter_n2), .ZN(
        extimating_unit_CU_adapter_ADD3_VALID_delay_2_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_VALID_delay_2_Q_int_reg ( .D(
        extimating_unit_CU_adapter_ADD3_VALID_int[1]), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_VALID_delay_2_n1), .Q(
        extimating_unit_CU_adapter_ADD3_VALID_int[2]) );
  INV_X1 extimating_unit_CU_adapter_ADD3_VALID_delay_3_U3 ( .A(
        extimating_unit_CU_adapter_n2), .ZN(
        extimating_unit_CU_adapter_ADD3_VALID_delay_3_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_VALID_delay_3_Q_int_reg ( .D(
        extimating_unit_CU_adapter_ADD3_VALID_int[2]), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_VALID_delay_3_n1), .Q(
        extimating_unit_CU_adapter_ADD3_VALID_int[3]) );
  INV_X1 extimating_unit_CU_adapter_ADD3_VALID_delay_4_U3 ( .A(
        extimating_unit_CU_adapter_n2), .ZN(
        extimating_unit_CU_adapter_ADD3_VALID_delay_4_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_VALID_delay_4_Q_int_reg ( .D(
        extimating_unit_CU_adapter_ADD3_VALID_int[3]), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_VALID_delay_4_n1), .Q(
        extimating_unit_CU_adapter_ADD3_VALID_int[4]) );
  INV_X1 extimating_unit_CU_adapter_ADD3_VALID_delay_5_U3 ( .A(
        extimating_unit_CU_adapter_n2), .ZN(
        extimating_unit_CU_adapter_ADD3_VALID_delay_5_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_VALID_delay_5_Q_int_reg ( .D(
        extimating_unit_CU_adapter_ADD3_VALID_int[4]), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_VALID_delay_5_n1), .Q(ADD3_VALID) );
  INV_X1 extimating_unit_CU_adapter_incrY_delay_1_U3 ( .A(
        extimating_unit_CU_adapter_n2), .ZN(
        extimating_unit_CU_adapter_incrY_delay_1_n1) );
  DFFR_X1 extimating_unit_CU_adapter_incrY_delay_1_Q_int_reg ( .D(ADD3_VALID), 
        .CK(clk), .RN(extimating_unit_CU_adapter_incrY_delay_1_n1), .Q(
        extimating_unit_CU_adapter_incrY_int[1]) );
  INV_X1 extimating_unit_CU_adapter_incrY_delay_2_U3 ( .A(
        extimating_unit_CU_adapter_n2), .ZN(
        extimating_unit_CU_adapter_incrY_delay_2_n1) );
  DFFR_X1 extimating_unit_CU_adapter_incrY_delay_2_Q_int_reg ( .D(
        extimating_unit_CU_adapter_incrY_int[1]), .CK(clk), .RN(
        extimating_unit_CU_adapter_incrY_delay_2_n1), .Q(
        extimating_unit_CU_adapter_incrY_int[2]) );
  INV_X1 extimating_unit_CU_adapter_incrY_delay_3_U3 ( .A(
        extimating_unit_CU_adapter_n3), .ZN(
        extimating_unit_CU_adapter_incrY_delay_3_n1) );
  DFFR_X1 extimating_unit_CU_adapter_incrY_delay_3_Q_int_reg ( .D(
        extimating_unit_CU_adapter_incrY_int[2]), .CK(clk), .RN(
        extimating_unit_CU_adapter_incrY_delay_3_n1), .Q(incrY) );
  INV_X1 extimating_unit_CU_adapter_MEM_RE_delay_1_U3 ( .A(
        extimating_unit_CU_adapter_n3), .ZN(
        extimating_unit_CU_adapter_MEM_RE_delay_1_n1) );
  DFFR_X1 extimating_unit_CU_adapter_MEM_RE_delay_1_Q_int_reg ( .D(incrY), 
        .CK(clk), .RN(extimating_unit_CU_adapter_MEM_RE_delay_1_n1), .Q(MEM_RE) );
  INV_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_1_U3 ( .A(
        extimating_unit_CU_adapter_n3), .ZN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_1_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_1_Q_int_reg ( .D(
        ADD3_MVin_LE_nSET), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_1_n1), .Q(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[1]) );
  INV_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_2_U3 ( .A(
        extimating_unit_CU_adapter_n3), .ZN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_2_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_2_Q_int_reg ( .D(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[1]), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_2_n1), .Q(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[2]) );
  INV_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_3_U3 ( .A(
        extimating_unit_CU_adapter_n3), .ZN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_3_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_3_Q_int_reg ( .D(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[2]), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_3_n1), .Q(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[3]) );
  INV_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_4_U3 ( .A(
        extimating_unit_CU_adapter_n3), .ZN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_4_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_4_Q_int_reg ( .D(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[3]), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_4_n1), .Q(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[4]) );
  INV_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_5_U3 ( .A(
        extimating_unit_CU_adapter_n3), .ZN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_5_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_5_Q_int_reg ( .D(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[4]), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_5_n1), .Q(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[5]) );
  INV_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_6_U3 ( .A(
        extimating_unit_CU_adapter_n3), .ZN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_6_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_6_Q_int_reg ( .D(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[5]), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_6_n1), .Q(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[6]) );
  INV_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_7_U3 ( .A(
        extimating_unit_CU_adapter_n3), .ZN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_7_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_7_Q_int_reg ( .D(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[6]), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_7_n1), .Q(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[7]) );
  INV_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_8_U3 ( .A(
        extimating_unit_CU_adapter_n3), .ZN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_8_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_8_Q_int_reg ( .D(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[7]), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_8_n1), .Q(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[8]) );
  INV_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_9_U3 ( .A(
        extimating_unit_CU_adapter_n3), .ZN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_9_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_9_Q_int_reg ( .D(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[8]), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_delay_9_n1), .Q(
        extimating_unit_CU_adapter_ADD3_MVin_LE_nSET_int[9]) );
  INV_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_register_U3 ( .A(
        extimating_unit_CU_adapter_ADD3_MVin_LE_fRESET_half_delayed), .ZN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_register_n1) );
  DFFR_X1 extimating_unit_CU_adapter_ADD3_MVin_LE_register_Q_int_reg ( .D(
        ADD3_MVin_LE), .CK(clk), .RN(
        extimating_unit_CU_adapter_ADD3_MVin_LE_register_n1), .Q(
        extimating_unit_CU_adapter_A3MVin_LE_samp) );
  INV_X1 extimating_unit_CU_adapter_LE_ab_delay_1_U3 ( .A(
        extimating_unit_CU_adapter_n3), .ZN(
        extimating_unit_CU_adapter_LE_ab_delay_1_n1) );
  DFFR_X1 extimating_unit_CU_adapter_LE_ab_delay_1_Q_int_reg ( .D(
        extimating_unit_LE_ab_CU_int), .CK(clk), .RN(
        extimating_unit_CU_adapter_LE_ab_delay_1_n1), .Q(
        extimating_unit_CU_adapter_LE_ab_int[1]) );
  INV_X1 extimating_unit_CU_adapter_LE_ab_delay_2_U3 ( .A(
        extimating_unit_CU_adapter_n4), .ZN(
        extimating_unit_CU_adapter_LE_ab_delay_2_n1) );
  DFFR_X1 extimating_unit_CU_adapter_LE_ab_delay_2_Q_int_reg ( .D(
        extimating_unit_CU_adapter_LE_ab_int[1]), .CK(clk), .RN(
        extimating_unit_CU_adapter_LE_ab_delay_2_n1), .Q(
        extimating_unit_CU_adapter_LE_ab_int[2]) );
  INV_X1 extimating_unit_CU_adapter_LE_ab_delay_3_U3 ( .A(
        extimating_unit_CU_adapter_n4), .ZN(
        extimating_unit_CU_adapter_LE_ab_delay_3_n1) );
  DFFR_X1 extimating_unit_CU_adapter_LE_ab_delay_3_Q_int_reg ( .D(
        extimating_unit_CU_adapter_LE_ab_int[2]), .CK(clk), .RN(
        extimating_unit_CU_adapter_LE_ab_delay_3_n1), .Q(
        extimating_unit_CU_adapter_LE_ab_int[3]) );
  INV_X1 extimating_unit_CU_adapter_LE_ab_delay_4_U3 ( .A(
        extimating_unit_CU_adapter_n4), .ZN(
        extimating_unit_CU_adapter_LE_ab_delay_4_n1) );
  DFFR_X1 extimating_unit_CU_adapter_LE_ab_delay_4_Q_int_reg ( .D(
        extimating_unit_CU_adapter_LE_ab_int[3]), .CK(clk), .RN(
        extimating_unit_CU_adapter_LE_ab_delay_4_n1), .Q(LE_ab) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_1_U3 ( .A(
        extimating_unit_CU_adapter_n4), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_1_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_1_Q_int_reg ( .D(
        extimating_unit_SAD_tmp_RST_CU_int), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_1_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[1]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_2_U3 ( .A(
        extimating_unit_CU_adapter_n4), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_2_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_2_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[1]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_2_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[2]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_3_U3 ( .A(
        extimating_unit_CU_adapter_n4), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_3_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_3_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[2]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_3_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[3]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_4_U3 ( .A(
        extimating_unit_CU_adapter_n4), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_4_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_4_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[3]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_4_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[4]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_5_U3 ( .A(
        extimating_unit_CU_adapter_n4), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_5_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_5_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[4]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_5_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[5]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_6_U3 ( .A(
        extimating_unit_CU_adapter_n4), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_6_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_6_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[5]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_6_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[6]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_7_U3 ( .A(
        extimating_unit_CU_adapter_n4), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_7_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_7_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[6]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_7_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[7]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_8_U3 ( .A(
        extimating_unit_CU_adapter_n4), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_8_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_8_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[7]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_8_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[8]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_9_U3 ( .A(
        extimating_unit_CU_adapter_n4), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_9_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_9_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[8]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_9_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[9]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_10_U3 ( .A(
        extimating_unit_CU_adapter_n5), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_10_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_10_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[9]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_10_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[10]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_11_U3 ( .A(
        extimating_unit_CU_adapter_n5), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_11_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_11_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[10]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_11_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[11]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_12_U3 ( .A(
        extimating_unit_CU_adapter_n5), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_12_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_12_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[11]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_12_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[12]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_13_U3 ( .A(
        extimating_unit_CU_adapter_n5), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_13_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_13_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[12]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_13_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[13]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_14_U3 ( .A(
        extimating_unit_CU_adapter_n5), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_14_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_14_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[13]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_14_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[14]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_15_U3 ( .A(
        extimating_unit_CU_adapter_n5), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_15_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_15_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[14]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_15_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[15]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_16_U3 ( .A(
        extimating_unit_CU_adapter_n5), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_16_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_16_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[15]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_16_n1), .Q(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[16]) );
  INV_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_17_U3 ( .A(
        extimating_unit_CU_adapter_n5), .ZN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_17_n1) );
  DFFR_X1 extimating_unit_CU_adapter_SAD_tmp_RST_delay_17_Q_int_reg ( .D(
        extimating_unit_CU_adapter_SAD_tmp_RST_int[16]), .CK(clk), .RN(
        extimating_unit_CU_adapter_SAD_tmp_RST_delay_17_n1), .Q(SAD_tmp_RST)
         );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_1_U3 ( .A(
        extimating_unit_CU_adapter_n5), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_1_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_1_Q_int_reg ( .D(
        INTER_DATA_VALID_RESET), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_1_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[1]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_2_U3 ( .A(
        extimating_unit_CU_adapter_n5), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_2_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_2_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[1]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_2_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[2]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_3_U3 ( .A(
        extimating_unit_CU_adapter_n5), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_3_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_3_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[2]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_3_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[3]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_4_U3 ( .A(
        extimating_unit_CU_adapter_n5), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_4_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_4_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[3]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_4_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[4]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_5_U3 ( .A(
        extimating_unit_CU_adapter_n6), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_5_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_5_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[4]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_5_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[5]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_6_U3 ( .A(
        extimating_unit_CU_adapter_n6), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_6_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_6_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[5]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_6_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[6]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_7_U3 ( .A(
        extimating_unit_CU_adapter_n6), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_7_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_7_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[6]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_7_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[7]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_8_U3 ( .A(
        extimating_unit_CU_adapter_n6), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_8_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_8_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[7]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_8_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[8]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_9_U3 ( .A(
        extimating_unit_CU_adapter_n6), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_9_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_9_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[8]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_9_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[9]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_10_U3 ( .A(
        extimating_unit_CU_adapter_n6), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_10_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_10_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[9]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_10_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[10]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_11_U3 ( .A(
        extimating_unit_CU_adapter_n6), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_11_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_11_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[10]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_11_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[11]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_12_U3 ( .A(
        extimating_unit_CU_adapter_n6), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_12_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_12_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[11]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_12_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[12]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_13_U3 ( .A(
        extimating_unit_CU_adapter_n6), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_13_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_13_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[12]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_13_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[13]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_14_U3 ( .A(
        extimating_unit_CU_adapter_n6), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_14_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_14_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[13]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_14_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[14]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_15_U3 ( .A(
        extimating_unit_CU_adapter_n6), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_15_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_15_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[14]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_15_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[15]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_16_U3 ( .A(
        extimating_unit_CU_adapter_n6), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_16_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_16_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[15]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_16_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[16]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_17_U3 ( .A(
        extimating_unit_CU_adapter_n9), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_17_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_17_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[16]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_17_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[17]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_18_U3 ( .A(
        extimating_unit_CU_adapter_n9), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_18_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_18_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[17]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_18_n1), .Q(
        extimating_unit_CU_adapter_Comp_EN_int[18]) );
  INV_X1 extimating_unit_CU_adapter_Comp_EN_delay_19_U3 ( .A(
        extimating_unit_CU_adapter_n9), .ZN(
        extimating_unit_CU_adapter_Comp_EN_delay_19_n1) );
  DFFR_X1 extimating_unit_CU_adapter_Comp_EN_delay_19_Q_int_reg ( .D(
        extimating_unit_CU_adapter_Comp_EN_int[18]), .CK(clk), .RN(
        extimating_unit_CU_adapter_Comp_EN_delay_19_n1), .Q(eComp_EN) );
  NAND2_X1 extimating_unit_Results_calculator_U153 ( .A1(
        extimating_unit_MV2_out_int[21]), .A2(
        extimating_unit_Results_calculator_n209), .ZN(
        extimating_unit_Results_calculator_n66) );
  OAI21_X1 extimating_unit_Results_calculator_U152 ( .B1(
        extimating_unit_Results_calculator_n132), .B2(
        extimating_unit_Results_calculator_n217), .A(
        extimating_unit_Results_calculator_n66), .ZN(
        extimating_unit_Results_calculator_n199) );
  NAND2_X1 extimating_unit_Results_calculator_U151 ( .A1(
        extimating_unit_MV2_out_int[20]), .A2(
        extimating_unit_Results_calculator_n207), .ZN(
        extimating_unit_Results_calculator_n65) );
  OAI21_X1 extimating_unit_Results_calculator_U150 ( .B1(
        extimating_unit_Results_calculator_n131), .B2(
        extimating_unit_Results_calculator_n217), .A(
        extimating_unit_Results_calculator_n65), .ZN(
        extimating_unit_Results_calculator_n197) );
  NAND2_X1 extimating_unit_Results_calculator_U149 ( .A1(
        extimating_unit_MV2_out_int[19]), .A2(
        extimating_unit_Results_calculator_n207), .ZN(
        extimating_unit_Results_calculator_n64) );
  OAI21_X1 extimating_unit_Results_calculator_U148 ( .B1(
        extimating_unit_Results_calculator_n130), .B2(
        extimating_unit_Results_calculator_n217), .A(
        extimating_unit_Results_calculator_n64), .ZN(
        extimating_unit_Results_calculator_n196) );
  NAND2_X1 extimating_unit_Results_calculator_U147 ( .A1(
        extimating_unit_MV2_out_int[18]), .A2(
        extimating_unit_Results_calculator_n207), .ZN(
        extimating_unit_Results_calculator_n63) );
  OAI21_X1 extimating_unit_Results_calculator_U146 ( .B1(
        extimating_unit_Results_calculator_n129), .B2(
        extimating_unit_Results_calculator_n217), .A(
        extimating_unit_Results_calculator_n63), .ZN(
        extimating_unit_Results_calculator_n195) );
  NAND2_X1 extimating_unit_Results_calculator_U145 ( .A1(
        extimating_unit_MV2_out_int[17]), .A2(
        extimating_unit_Results_calculator_n207), .ZN(
        extimating_unit_Results_calculator_n62) );
  OAI21_X1 extimating_unit_Results_calculator_U144 ( .B1(
        extimating_unit_Results_calculator_n128), .B2(
        extimating_unit_Results_calculator_n217), .A(
        extimating_unit_Results_calculator_n62), .ZN(
        extimating_unit_Results_calculator_n194) );
  NAND2_X1 extimating_unit_Results_calculator_U143 ( .A1(
        extimating_unit_MV2_out_int[16]), .A2(
        extimating_unit_Results_calculator_n207), .ZN(
        extimating_unit_Results_calculator_n61) );
  OAI21_X1 extimating_unit_Results_calculator_U142 ( .B1(
        extimating_unit_Results_calculator_n127), .B2(
        extimating_unit_Results_calculator_n217), .A(
        extimating_unit_Results_calculator_n61), .ZN(
        extimating_unit_Results_calculator_n193) );
  NAND2_X1 extimating_unit_Results_calculator_U141 ( .A1(
        extimating_unit_MV2_out_int[15]), .A2(
        extimating_unit_Results_calculator_n207), .ZN(
        extimating_unit_Results_calculator_n60) );
  OAI21_X1 extimating_unit_Results_calculator_U140 ( .B1(
        extimating_unit_Results_calculator_n126), .B2(
        extimating_unit_Results_calculator_n216), .A(
        extimating_unit_Results_calculator_n60), .ZN(
        extimating_unit_Results_calculator_n192) );
  NAND2_X1 extimating_unit_Results_calculator_U139 ( .A1(
        extimating_unit_MV2_out_int[14]), .A2(
        extimating_unit_Results_calculator_n207), .ZN(
        extimating_unit_Results_calculator_n59) );
  OAI21_X1 extimating_unit_Results_calculator_U138 ( .B1(
        extimating_unit_Results_calculator_n125), .B2(
        extimating_unit_Results_calculator_n217), .A(
        extimating_unit_Results_calculator_n59), .ZN(
        extimating_unit_Results_calculator_n191) );
  NAND2_X1 extimating_unit_Results_calculator_U137 ( .A1(
        extimating_unit_MV2_out_int[13]), .A2(
        extimating_unit_Results_calculator_n207), .ZN(
        extimating_unit_Results_calculator_n58) );
  OAI21_X1 extimating_unit_Results_calculator_U135 ( .B1(
        extimating_unit_Results_calculator_n124), .B2(
        extimating_unit_Results_calculator_n216), .A(
        extimating_unit_Results_calculator_n58), .ZN(
        extimating_unit_Results_calculator_n190) );
  NAND2_X1 extimating_unit_Results_calculator_U134 ( .A1(
        extimating_unit_MV2_out_int[12]), .A2(
        extimating_unit_Results_calculator_n207), .ZN(
        extimating_unit_Results_calculator_n57) );
  OAI21_X1 extimating_unit_Results_calculator_U133 ( .B1(
        extimating_unit_Results_calculator_n123), .B2(
        extimating_unit_Results_calculator_n216), .A(
        extimating_unit_Results_calculator_n57), .ZN(
        extimating_unit_Results_calculator_n189) );
  NAND2_X1 extimating_unit_Results_calculator_U132 ( .A1(
        extimating_unit_MV2_out_int[11]), .A2(
        extimating_unit_Results_calculator_n207), .ZN(
        extimating_unit_Results_calculator_n56) );
  OAI21_X1 extimating_unit_Results_calculator_U131 ( .B1(
        extimating_unit_Results_calculator_n122), .B2(
        extimating_unit_Results_calculator_n216), .A(
        extimating_unit_Results_calculator_n56), .ZN(
        extimating_unit_Results_calculator_n188) );
  NAND2_X1 extimating_unit_Results_calculator_U130 ( .A1(
        extimating_unit_MV2_out_int[10]), .A2(
        extimating_unit_Results_calculator_n207), .ZN(
        extimating_unit_Results_calculator_n55) );
  OAI21_X1 extimating_unit_Results_calculator_U129 ( .B1(
        extimating_unit_Results_calculator_n121), .B2(
        extimating_unit_Results_calculator_n216), .A(
        extimating_unit_Results_calculator_n55), .ZN(
        extimating_unit_Results_calculator_n187) );
  NAND2_X1 extimating_unit_Results_calculator_U128 ( .A1(
        extimating_unit_MV2_out_int[9]), .A2(
        extimating_unit_Results_calculator_n207), .ZN(
        extimating_unit_Results_calculator_n54) );
  OAI21_X1 extimating_unit_Results_calculator_U127 ( .B1(
        extimating_unit_Results_calculator_n120), .B2(
        extimating_unit_Results_calculator_n216), .A(
        extimating_unit_Results_calculator_n54), .ZN(
        extimating_unit_Results_calculator_n186) );
  NAND2_X1 extimating_unit_Results_calculator_U126 ( .A1(
        extimating_unit_MV2_out_int[8]), .A2(
        extimating_unit_Results_calculator_n208), .ZN(
        extimating_unit_Results_calculator_n53) );
  OAI21_X1 extimating_unit_Results_calculator_U125 ( .B1(
        extimating_unit_Results_calculator_n119), .B2(
        extimating_unit_Results_calculator_n216), .A(
        extimating_unit_Results_calculator_n53), .ZN(
        extimating_unit_Results_calculator_n185) );
  NAND2_X1 extimating_unit_Results_calculator_U124 ( .A1(
        extimating_unit_MV2_out_int[7]), .A2(
        extimating_unit_Results_calculator_n208), .ZN(
        extimating_unit_Results_calculator_n52) );
  OAI21_X1 extimating_unit_Results_calculator_U123 ( .B1(
        extimating_unit_Results_calculator_n118), .B2(
        extimating_unit_Results_calculator_n215), .A(
        extimating_unit_Results_calculator_n52), .ZN(
        extimating_unit_Results_calculator_n184) );
  NAND2_X1 extimating_unit_Results_calculator_U122 ( .A1(
        extimating_unit_MV2_out_int[6]), .A2(
        extimating_unit_Results_calculator_n208), .ZN(
        extimating_unit_Results_calculator_n51) );
  OAI21_X1 extimating_unit_Results_calculator_U121 ( .B1(
        extimating_unit_Results_calculator_n117), .B2(
        extimating_unit_Results_calculator_n215), .A(
        extimating_unit_Results_calculator_n51), .ZN(
        extimating_unit_Results_calculator_n183) );
  NAND2_X1 extimating_unit_Results_calculator_U120 ( .A1(
        extimating_unit_MV2_out_int[5]), .A2(
        extimating_unit_Results_calculator_n208), .ZN(
        extimating_unit_Results_calculator_n50) );
  OAI21_X1 extimating_unit_Results_calculator_U119 ( .B1(
        extimating_unit_Results_calculator_n116), .B2(
        extimating_unit_Results_calculator_n216), .A(
        extimating_unit_Results_calculator_n50), .ZN(
        extimating_unit_Results_calculator_n182) );
  NAND2_X1 extimating_unit_Results_calculator_U118 ( .A1(
        extimating_unit_MV2_out_int[4]), .A2(
        extimating_unit_Results_calculator_n208), .ZN(
        extimating_unit_Results_calculator_n49) );
  OAI21_X1 extimating_unit_Results_calculator_U117 ( .B1(
        extimating_unit_Results_calculator_n115), .B2(
        extimating_unit_Results_calculator_n215), .A(
        extimating_unit_Results_calculator_n49), .ZN(
        extimating_unit_Results_calculator_n181) );
  NAND2_X1 extimating_unit_Results_calculator_U116 ( .A1(
        extimating_unit_MV2_out_int[3]), .A2(
        extimating_unit_Results_calculator_n208), .ZN(
        extimating_unit_Results_calculator_n48) );
  OAI21_X1 extimating_unit_Results_calculator_U115 ( .B1(
        extimating_unit_Results_calculator_n114), .B2(
        extimating_unit_Results_calculator_n215), .A(
        extimating_unit_Results_calculator_n48), .ZN(
        extimating_unit_Results_calculator_n180) );
  NAND2_X1 extimating_unit_Results_calculator_U114 ( .A1(
        extimating_unit_MV2_out_int[2]), .A2(
        extimating_unit_Results_calculator_n208), .ZN(
        extimating_unit_Results_calculator_n47) );
  OAI21_X1 extimating_unit_Results_calculator_U113 ( .B1(
        extimating_unit_Results_calculator_n113), .B2(
        extimating_unit_Results_calculator_n215), .A(
        extimating_unit_Results_calculator_n47), .ZN(
        extimating_unit_Results_calculator_n179) );
  NAND2_X1 extimating_unit_Results_calculator_U112 ( .A1(
        extimating_unit_MV2_out_int[1]), .A2(
        extimating_unit_Results_calculator_n208), .ZN(
        extimating_unit_Results_calculator_n46) );
  OAI21_X1 extimating_unit_Results_calculator_U111 ( .B1(
        extimating_unit_Results_calculator_n112), .B2(
        extimating_unit_Results_calculator_n215), .A(
        extimating_unit_Results_calculator_n46), .ZN(
        extimating_unit_Results_calculator_n178) );
  NAND2_X1 extimating_unit_Results_calculator_U110 ( .A1(
        extimating_unit_MV2_out_int[0]), .A2(
        extimating_unit_Results_calculator_n208), .ZN(
        extimating_unit_Results_calculator_n45) );
  OAI21_X1 extimating_unit_Results_calculator_U109 ( .B1(
        extimating_unit_Results_calculator_n111), .B2(
        extimating_unit_Results_calculator_n214), .A(
        extimating_unit_Results_calculator_n45), .ZN(
        extimating_unit_Results_calculator_n177) );
  NAND2_X1 extimating_unit_Results_calculator_U108 ( .A1(
        extimating_unit_MV0_out_int[21]), .A2(
        extimating_unit_Results_calculator_n208), .ZN(
        extimating_unit_Results_calculator_n44) );
  OAI21_X1 extimating_unit_Results_calculator_U107 ( .B1(
        extimating_unit_Results_calculator_n110), .B2(
        extimating_unit_Results_calculator_n215), .A(
        extimating_unit_Results_calculator_n44), .ZN(
        extimating_unit_Results_calculator_n176) );
  NAND2_X1 extimating_unit_Results_calculator_U106 ( .A1(
        extimating_unit_MV0_out_int[20]), .A2(
        extimating_unit_Results_calculator_n208), .ZN(
        extimating_unit_Results_calculator_n43) );
  OAI21_X1 extimating_unit_Results_calculator_U105 ( .B1(
        extimating_unit_Results_calculator_n109), .B2(
        extimating_unit_Results_calculator_n214), .A(
        extimating_unit_Results_calculator_n43), .ZN(
        extimating_unit_Results_calculator_n175) );
  NAND2_X1 extimating_unit_Results_calculator_U104 ( .A1(
        extimating_unit_MV0_out_int[19]), .A2(
        extimating_unit_Results_calculator_n208), .ZN(
        extimating_unit_Results_calculator_n42) );
  OAI21_X1 extimating_unit_Results_calculator_U103 ( .B1(
        extimating_unit_Results_calculator_n108), .B2(
        extimating_unit_Results_calculator_n214), .A(
        extimating_unit_Results_calculator_n42), .ZN(
        extimating_unit_Results_calculator_n174) );
  NAND2_X1 extimating_unit_Results_calculator_U102 ( .A1(
        extimating_unit_MV0_out_int[18]), .A2(
        extimating_unit_Results_calculator_n209), .ZN(
        extimating_unit_Results_calculator_n41) );
  OAI21_X1 extimating_unit_Results_calculator_U101 ( .B1(
        extimating_unit_Results_calculator_n107), .B2(
        extimating_unit_Results_calculator_n214), .A(
        extimating_unit_Results_calculator_n41), .ZN(
        extimating_unit_Results_calculator_n173) );
  NAND2_X1 extimating_unit_Results_calculator_U100 ( .A1(
        extimating_unit_MV0_out_int[17]), .A2(
        extimating_unit_Results_calculator_n209), .ZN(
        extimating_unit_Results_calculator_n40) );
  OAI21_X1 extimating_unit_Results_calculator_U99 ( .B1(
        extimating_unit_Results_calculator_n106), .B2(
        extimating_unit_Results_calculator_n214), .A(
        extimating_unit_Results_calculator_n40), .ZN(
        extimating_unit_Results_calculator_n172) );
  NAND2_X1 extimating_unit_Results_calculator_U98 ( .A1(
        extimating_unit_MV0_out_int[16]), .A2(
        extimating_unit_Results_calculator_n209), .ZN(
        extimating_unit_Results_calculator_n39) );
  OAI21_X1 extimating_unit_Results_calculator_U97 ( .B1(
        extimating_unit_Results_calculator_n105), .B2(
        extimating_unit_Results_calculator_n214), .A(
        extimating_unit_Results_calculator_n39), .ZN(
        extimating_unit_Results_calculator_n171) );
  NAND2_X1 extimating_unit_Results_calculator_U96 ( .A1(
        extimating_unit_MV0_out_int[15]), .A2(
        extimating_unit_Results_calculator_n209), .ZN(
        extimating_unit_Results_calculator_n38) );
  OAI21_X1 extimating_unit_Results_calculator_U95 ( .B1(
        extimating_unit_Results_calculator_n104), .B2(
        extimating_unit_Results_calculator_n214), .A(
        extimating_unit_Results_calculator_n38), .ZN(
        extimating_unit_Results_calculator_n170) );
  NAND2_X1 extimating_unit_Results_calculator_U94 ( .A1(
        extimating_unit_MV0_out_int[14]), .A2(
        extimating_unit_Results_calculator_n209), .ZN(
        extimating_unit_Results_calculator_n37) );
  OAI21_X1 extimating_unit_Results_calculator_U93 ( .B1(
        extimating_unit_Results_calculator_n103), .B2(
        extimating_unit_Results_calculator_n213), .A(
        extimating_unit_Results_calculator_n37), .ZN(
        extimating_unit_Results_calculator_n169) );
  NAND2_X1 extimating_unit_Results_calculator_U92 ( .A1(
        extimating_unit_MV0_out_int[13]), .A2(
        extimating_unit_Results_calculator_n209), .ZN(
        extimating_unit_Results_calculator_n36) );
  OAI21_X1 extimating_unit_Results_calculator_U91 ( .B1(
        extimating_unit_Results_calculator_n102), .B2(
        extimating_unit_Results_calculator_n213), .A(
        extimating_unit_Results_calculator_n36), .ZN(
        extimating_unit_Results_calculator_n168) );
  NAND2_X1 extimating_unit_Results_calculator_U90 ( .A1(
        extimating_unit_MV0_out_int[12]), .A2(
        extimating_unit_Results_calculator_n209), .ZN(
        extimating_unit_Results_calculator_n35) );
  OAI21_X1 extimating_unit_Results_calculator_U89 ( .B1(
        extimating_unit_Results_calculator_n101), .B2(
        extimating_unit_Results_calculator_n214), .A(
        extimating_unit_Results_calculator_n35), .ZN(
        extimating_unit_Results_calculator_n167) );
  NAND2_X1 extimating_unit_Results_calculator_U88 ( .A1(
        extimating_unit_MV0_out_int[11]), .A2(
        extimating_unit_Results_calculator_n209), .ZN(
        extimating_unit_Results_calculator_n34) );
  OAI21_X1 extimating_unit_Results_calculator_U87 ( .B1(
        extimating_unit_Results_calculator_n100), .B2(
        extimating_unit_Results_calculator_n213), .A(
        extimating_unit_Results_calculator_n34), .ZN(
        extimating_unit_Results_calculator_n166) );
  NAND2_X1 extimating_unit_Results_calculator_U86 ( .A1(
        extimating_unit_MV0_out_int[10]), .A2(
        extimating_unit_Results_calculator_n210), .ZN(
        extimating_unit_Results_calculator_n33) );
  OAI21_X1 extimating_unit_Results_calculator_U85 ( .B1(
        extimating_unit_Results_calculator_n99), .B2(
        extimating_unit_Results_calculator_n213), .A(
        extimating_unit_Results_calculator_n33), .ZN(
        extimating_unit_Results_calculator_n165) );
  NAND2_X1 extimating_unit_Results_calculator_U84 ( .A1(
        extimating_unit_MV0_out_int[9]), .A2(
        extimating_unit_Results_calculator_n209), .ZN(
        extimating_unit_Results_calculator_n32) );
  OAI21_X1 extimating_unit_Results_calculator_U83 ( .B1(
        extimating_unit_Results_calculator_n98), .B2(
        extimating_unit_Results_calculator_n214), .A(
        extimating_unit_Results_calculator_n32), .ZN(
        extimating_unit_Results_calculator_n164) );
  NAND2_X1 extimating_unit_Results_calculator_U82 ( .A1(
        extimating_unit_MV0_out_int[8]), .A2(
        extimating_unit_Results_calculator_n209), .ZN(
        extimating_unit_Results_calculator_n31) );
  OAI21_X1 extimating_unit_Results_calculator_U81 ( .B1(
        extimating_unit_Results_calculator_n97), .B2(
        extimating_unit_Results_calculator_n212), .A(
        extimating_unit_Results_calculator_n31), .ZN(
        extimating_unit_Results_calculator_n163) );
  NAND2_X1 extimating_unit_Results_calculator_U80 ( .A1(
        extimating_unit_MV0_out_int[7]), .A2(
        extimating_unit_Results_calculator_n209), .ZN(
        extimating_unit_Results_calculator_n30) );
  OAI21_X1 extimating_unit_Results_calculator_U79 ( .B1(
        extimating_unit_Results_calculator_n96), .B2(
        extimating_unit_Results_calculator_n212), .A(
        extimating_unit_Results_calculator_n30), .ZN(
        extimating_unit_Results_calculator_n162) );
  NAND2_X1 extimating_unit_Results_calculator_U78 ( .A1(
        extimating_unit_MV0_out_int[6]), .A2(
        extimating_unit_Results_calculator_n210), .ZN(
        extimating_unit_Results_calculator_n29) );
  OAI21_X1 extimating_unit_Results_calculator_U77 ( .B1(
        extimating_unit_Results_calculator_n95), .B2(
        extimating_unit_Results_calculator_n213), .A(
        extimating_unit_Results_calculator_n29), .ZN(
        extimating_unit_Results_calculator_n161) );
  NAND2_X1 extimating_unit_Results_calculator_U76 ( .A1(
        extimating_unit_MV0_out_int[5]), .A2(
        extimating_unit_Results_calculator_n210), .ZN(
        extimating_unit_Results_calculator_n28) );
  OAI21_X1 extimating_unit_Results_calculator_U75 ( .B1(
        extimating_unit_Results_calculator_n94), .B2(
        extimating_unit_Results_calculator_n212), .A(
        extimating_unit_Results_calculator_n28), .ZN(
        extimating_unit_Results_calculator_n160) );
  NAND2_X1 extimating_unit_Results_calculator_U74 ( .A1(
        extimating_unit_MV0_out_int[4]), .A2(
        extimating_unit_Results_calculator_n210), .ZN(
        extimating_unit_Results_calculator_n27) );
  OAI21_X1 extimating_unit_Results_calculator_U73 ( .B1(
        extimating_unit_Results_calculator_n93), .B2(
        extimating_unit_Results_calculator_n212), .A(
        extimating_unit_Results_calculator_n27), .ZN(
        extimating_unit_Results_calculator_n159) );
  NAND2_X1 extimating_unit_Results_calculator_U72 ( .A1(
        extimating_unit_MV0_out_int[3]), .A2(
        extimating_unit_Results_calculator_n210), .ZN(
        extimating_unit_Results_calculator_n26) );
  OAI21_X1 extimating_unit_Results_calculator_U71 ( .B1(
        extimating_unit_Results_calculator_n92), .B2(
        extimating_unit_Results_calculator_n213), .A(
        extimating_unit_Results_calculator_n26), .ZN(
        extimating_unit_Results_calculator_n158) );
  NAND2_X1 extimating_unit_Results_calculator_U70 ( .A1(
        extimating_unit_MV0_out_int[2]), .A2(
        extimating_unit_Results_calculator_n210), .ZN(
        extimating_unit_Results_calculator_n25) );
  OAI21_X1 extimating_unit_Results_calculator_U69 ( .B1(
        extimating_unit_Results_calculator_n91), .B2(
        extimating_unit_Results_calculator_n212), .A(
        extimating_unit_Results_calculator_n25), .ZN(
        extimating_unit_Results_calculator_n157) );
  NAND2_X1 extimating_unit_Results_calculator_U68 ( .A1(
        extimating_unit_MV0_out_int[1]), .A2(
        extimating_unit_Results_calculator_n210), .ZN(
        extimating_unit_Results_calculator_n24) );
  OAI21_X1 extimating_unit_Results_calculator_U67 ( .B1(
        extimating_unit_Results_calculator_n90), .B2(
        extimating_unit_Results_calculator_n212), .A(
        extimating_unit_Results_calculator_n24), .ZN(
        extimating_unit_Results_calculator_n156) );
  NAND2_X1 extimating_unit_Results_calculator_U66 ( .A1(
        extimating_unit_MV0_out_int[0]), .A2(
        extimating_unit_Results_calculator_n210), .ZN(
        extimating_unit_Results_calculator_n23) );
  OAI21_X1 extimating_unit_Results_calculator_U65 ( .B1(
        extimating_unit_Results_calculator_n89), .B2(
        extimating_unit_Results_calculator_n213), .A(
        extimating_unit_Results_calculator_n23), .ZN(
        extimating_unit_Results_calculator_n155) );
  NAND2_X1 extimating_unit_Results_calculator_U64 ( .A1(
        extimating_unit_MV1_out_int[21]), .A2(
        extimating_unit_Results_calculator_n210), .ZN(
        extimating_unit_Results_calculator_n22) );
  OAI21_X1 extimating_unit_Results_calculator_U63 ( .B1(
        extimating_unit_Results_calculator_n88), .B2(
        extimating_unit_Results_calculator_n213), .A(
        extimating_unit_Results_calculator_n22), .ZN(
        extimating_unit_Results_calculator_n154) );
  NAND2_X1 extimating_unit_Results_calculator_U62 ( .A1(
        extimating_unit_MV1_out_int[20]), .A2(
        extimating_unit_Results_calculator_n210), .ZN(
        extimating_unit_Results_calculator_n21) );
  OAI21_X1 extimating_unit_Results_calculator_U61 ( .B1(
        extimating_unit_Results_calculator_n87), .B2(
        extimating_unit_Results_calculator_n213), .A(
        extimating_unit_Results_calculator_n21), .ZN(
        extimating_unit_Results_calculator_n153) );
  NAND2_X1 extimating_unit_Results_calculator_U60 ( .A1(
        extimating_unit_MV1_out_int[19]), .A2(
        extimating_unit_Results_calculator_n210), .ZN(
        extimating_unit_Results_calculator_n20) );
  OAI21_X1 extimating_unit_Results_calculator_U59 ( .B1(
        extimating_unit_Results_calculator_n86), .B2(
        extimating_unit_Results_calculator_n212), .A(
        extimating_unit_Results_calculator_n20), .ZN(
        extimating_unit_Results_calculator_n152) );
  NAND2_X1 extimating_unit_Results_calculator_U58 ( .A1(
        extimating_unit_MV1_out_int[18]), .A2(
        extimating_unit_Results_calculator_n211), .ZN(
        extimating_unit_Results_calculator_n19) );
  OAI21_X1 extimating_unit_Results_calculator_U57 ( .B1(
        extimating_unit_Results_calculator_n85), .B2(
        extimating_unit_Results_calculator_n215), .A(
        extimating_unit_Results_calculator_n19), .ZN(
        extimating_unit_Results_calculator_n151) );
  NAND2_X1 extimating_unit_Results_calculator_U56 ( .A1(
        extimating_unit_MV1_out_int[17]), .A2(
        extimating_unit_Results_calculator_n211), .ZN(
        extimating_unit_Results_calculator_n18) );
  OAI21_X1 extimating_unit_Results_calculator_U55 ( .B1(
        extimating_unit_Results_calculator_n84), .B2(
        extimating_unit_Results_calculator_n213), .A(
        extimating_unit_Results_calculator_n18), .ZN(
        extimating_unit_Results_calculator_n150) );
  NAND2_X1 extimating_unit_Results_calculator_U54 ( .A1(
        extimating_unit_MV1_out_int[16]), .A2(
        extimating_unit_Results_calculator_n210), .ZN(
        extimating_unit_Results_calculator_n17) );
  OAI21_X1 extimating_unit_Results_calculator_U53 ( .B1(
        extimating_unit_Results_calculator_n83), .B2(
        extimating_unit_Results_calculator_n213), .A(
        extimating_unit_Results_calculator_n17), .ZN(
        extimating_unit_Results_calculator_n149) );
  NAND2_X1 extimating_unit_Results_calculator_U52 ( .A1(
        extimating_unit_MV1_out_int[15]), .A2(
        extimating_unit_Results_calculator_n211), .ZN(
        extimating_unit_Results_calculator_n16) );
  OAI21_X1 extimating_unit_Results_calculator_U51 ( .B1(
        extimating_unit_Results_calculator_n82), .B2(
        extimating_unit_Results_calculator_n214), .A(
        extimating_unit_Results_calculator_n16), .ZN(
        extimating_unit_Results_calculator_n148) );
  NAND2_X1 extimating_unit_Results_calculator_U50 ( .A1(
        extimating_unit_MV1_out_int[14]), .A2(
        extimating_unit_Results_calculator_n211), .ZN(
        extimating_unit_Results_calculator_n15) );
  OAI21_X1 extimating_unit_Results_calculator_U49 ( .B1(
        extimating_unit_Results_calculator_n81), .B2(
        extimating_unit_Results_calculator_n213), .A(
        extimating_unit_Results_calculator_n15), .ZN(
        extimating_unit_Results_calculator_n147) );
  NAND2_X1 extimating_unit_Results_calculator_U48 ( .A1(
        extimating_unit_MV1_out_int[13]), .A2(
        extimating_unit_Results_calculator_n211), .ZN(
        extimating_unit_Results_calculator_n14) );
  OAI21_X1 extimating_unit_Results_calculator_U47 ( .B1(
        extimating_unit_Results_calculator_n80), .B2(
        extimating_unit_Results_calculator_n214), .A(
        extimating_unit_Results_calculator_n14), .ZN(
        extimating_unit_Results_calculator_n146) );
  NAND2_X1 extimating_unit_Results_calculator_U46 ( .A1(
        extimating_unit_MV1_out_int[12]), .A2(
        extimating_unit_Results_calculator_n211), .ZN(
        extimating_unit_Results_calculator_n13) );
  OAI21_X1 extimating_unit_Results_calculator_U45 ( .B1(
        extimating_unit_Results_calculator_n79), .B2(
        extimating_unit_Results_calculator_n215), .A(
        extimating_unit_Results_calculator_n13), .ZN(
        extimating_unit_Results_calculator_n145) );
  NAND2_X1 extimating_unit_Results_calculator_U44 ( .A1(
        extimating_unit_MV1_out_int[11]), .A2(
        extimating_unit_Results_calculator_n211), .ZN(
        extimating_unit_Results_calculator_n12) );
  OAI21_X1 extimating_unit_Results_calculator_U43 ( .B1(
        extimating_unit_Results_calculator_n78), .B2(
        extimating_unit_Results_calculator_n214), .A(
        extimating_unit_Results_calculator_n12), .ZN(
        extimating_unit_Results_calculator_n144) );
  NAND2_X1 extimating_unit_Results_calculator_U42 ( .A1(
        extimating_unit_MV1_out_int[10]), .A2(
        extimating_unit_Results_calculator_n211), .ZN(
        extimating_unit_Results_calculator_n11) );
  OAI21_X1 extimating_unit_Results_calculator_U41 ( .B1(
        extimating_unit_Results_calculator_n77), .B2(
        extimating_unit_Results_calculator_n215), .A(
        extimating_unit_Results_calculator_n11), .ZN(
        extimating_unit_Results_calculator_n143) );
  NAND2_X1 extimating_unit_Results_calculator_U40 ( .A1(
        extimating_unit_MV1_out_int[9]), .A2(
        extimating_unit_Results_calculator_n211), .ZN(
        extimating_unit_Results_calculator_n10) );
  OAI21_X1 extimating_unit_Results_calculator_U39 ( .B1(
        extimating_unit_Results_calculator_n76), .B2(
        extimating_unit_Results_calculator_n216), .A(
        extimating_unit_Results_calculator_n10), .ZN(
        extimating_unit_Results_calculator_n142) );
  NAND2_X1 extimating_unit_Results_calculator_U38 ( .A1(
        extimating_unit_MV1_out_int[8]), .A2(
        extimating_unit_Results_calculator_n212), .ZN(
        extimating_unit_Results_calculator_n9) );
  OAI21_X1 extimating_unit_Results_calculator_U37 ( .B1(
        extimating_unit_Results_calculator_n75), .B2(
        extimating_unit_Results_calculator_n215), .A(
        extimating_unit_Results_calculator_n9), .ZN(
        extimating_unit_Results_calculator_n141) );
  NAND2_X1 extimating_unit_Results_calculator_U36 ( .A1(
        extimating_unit_MV1_out_int[7]), .A2(
        extimating_unit_Results_calculator_n211), .ZN(
        extimating_unit_Results_calculator_n8) );
  OAI21_X1 extimating_unit_Results_calculator_U35 ( .B1(
        extimating_unit_Results_calculator_n74), .B2(
        extimating_unit_Results_calculator_n215), .A(
        extimating_unit_Results_calculator_n8), .ZN(
        extimating_unit_Results_calculator_n140) );
  NAND2_X1 extimating_unit_Results_calculator_U34 ( .A1(
        extimating_unit_MV1_out_int[6]), .A2(
        extimating_unit_Results_calculator_n212), .ZN(
        extimating_unit_Results_calculator_n7) );
  OAI21_X1 extimating_unit_Results_calculator_U33 ( .B1(
        extimating_unit_Results_calculator_n73), .B2(
        extimating_unit_Results_calculator_n216), .A(
        extimating_unit_Results_calculator_n7), .ZN(
        extimating_unit_Results_calculator_n139) );
  NAND2_X1 extimating_unit_Results_calculator_U32 ( .A1(
        extimating_unit_MV1_out_int[5]), .A2(
        extimating_unit_Results_calculator_n212), .ZN(
        extimating_unit_Results_calculator_n6) );
  OAI21_X1 extimating_unit_Results_calculator_U31 ( .B1(
        extimating_unit_Results_calculator_n72), .B2(
        extimating_unit_Results_calculator_n216), .A(
        extimating_unit_Results_calculator_n6), .ZN(
        extimating_unit_Results_calculator_n138) );
  NAND2_X1 extimating_unit_Results_calculator_U30 ( .A1(
        extimating_unit_MV1_out_int[4]), .A2(
        extimating_unit_Results_calculator_n211), .ZN(
        extimating_unit_Results_calculator_n5) );
  OAI21_X1 extimating_unit_Results_calculator_U29 ( .B1(
        extimating_unit_Results_calculator_n71), .B2(
        extimating_unit_Results_calculator_n216), .A(
        extimating_unit_Results_calculator_n5), .ZN(
        extimating_unit_Results_calculator_n137) );
  NAND2_X1 extimating_unit_Results_calculator_U28 ( .A1(
        extimating_unit_MV1_out_int[3]), .A2(
        extimating_unit_Results_calculator_n212), .ZN(
        extimating_unit_Results_calculator_n4) );
  OAI21_X1 extimating_unit_Results_calculator_U27 ( .B1(
        extimating_unit_Results_calculator_n70), .B2(
        extimating_unit_Results_calculator_n217), .A(
        extimating_unit_Results_calculator_n4), .ZN(
        extimating_unit_Results_calculator_n136) );
  NAND2_X1 extimating_unit_Results_calculator_U26 ( .A1(
        extimating_unit_MV1_out_int[2]), .A2(
        extimating_unit_Results_calculator_n212), .ZN(
        extimating_unit_Results_calculator_n3) );
  OAI21_X1 extimating_unit_Results_calculator_U25 ( .B1(
        extimating_unit_Results_calculator_n69), .B2(
        extimating_unit_Results_calculator_n217), .A(
        extimating_unit_Results_calculator_n3), .ZN(
        extimating_unit_Results_calculator_n135) );
  NAND2_X1 extimating_unit_Results_calculator_U24 ( .A1(
        extimating_unit_MV1_out_int[1]), .A2(
        extimating_unit_Results_calculator_n211), .ZN(
        extimating_unit_Results_calculator_n2) );
  OAI21_X1 extimating_unit_Results_calculator_U23 ( .B1(
        extimating_unit_Results_calculator_n68), .B2(
        extimating_unit_Results_calculator_n217), .A(
        extimating_unit_Results_calculator_n2), .ZN(
        extimating_unit_Results_calculator_n134) );
  NAND2_X1 extimating_unit_Results_calculator_U22 ( .A1(
        extimating_unit_Results_calculator_n217), .A2(
        extimating_unit_MV1_out_int[0]), .ZN(
        extimating_unit_Results_calculator_n1) );
  OAI21_X1 extimating_unit_Results_calculator_U21 ( .B1(
        extimating_unit_Results_calculator_n67), .B2(
        extimating_unit_Results_calculator_n217), .A(
        extimating_unit_Results_calculator_n1), .ZN(
        extimating_unit_Results_calculator_n133) );
  AND2_X1 extimating_unit_Results_calculator_U20 ( .A1(
        extimating_unit_Results_calculator_ltmin), .A2(eComp_EN), .ZN(
        extimating_unit_Results_calculator_Found_best) );
  BUF_X1 extimating_unit_Results_calculator_U19 ( .A(extimating_unit_RST2_int), 
        .Z(extimating_unit_Results_calculator_n198) );
  BUF_X1 extimating_unit_Results_calculator_U18 ( .A(OUT_LE), .Z(
        extimating_unit_Results_calculator_n206) );
  BUF_X1 extimating_unit_Results_calculator_U17 ( .A(OUT_LE), .Z(
        extimating_unit_Results_calculator_n205) );
  BUF_X1 extimating_unit_Results_calculator_U16 ( .A(
        extimating_unit_Results_calculator_n198), .Z(
        extimating_unit_Results_calculator_n204) );
  BUF_X1 extimating_unit_Results_calculator_U15 ( .A(
        extimating_unit_Results_calculator_n198), .Z(
        extimating_unit_Results_calculator_n202) );
  BUF_X1 extimating_unit_Results_calculator_U14 ( .A(
        extimating_unit_Results_calculator_n198), .Z(
        extimating_unit_Results_calculator_n203) );
  BUF_X1 extimating_unit_Results_calculator_U13 ( .A(
        extimating_unit_Results_calculator_n206), .Z(
        extimating_unit_Results_calculator_n217) );
  BUF_X1 extimating_unit_Results_calculator_U12 ( .A(
        extimating_unit_Results_calculator_n206), .Z(
        extimating_unit_Results_calculator_n216) );
  BUF_X1 extimating_unit_Results_calculator_U11 ( .A(
        extimating_unit_Results_calculator_n206), .Z(
        extimating_unit_Results_calculator_n215) );
  BUF_X1 extimating_unit_Results_calculator_U10 ( .A(
        extimating_unit_Results_calculator_n206), .Z(
        extimating_unit_Results_calculator_n214) );
  BUF_X1 extimating_unit_Results_calculator_U9 ( .A(
        extimating_unit_Results_calculator_n206), .Z(
        extimating_unit_Results_calculator_n213) );
  BUF_X1 extimating_unit_Results_calculator_U8 ( .A(
        extimating_unit_Results_calculator_n205), .Z(
        extimating_unit_Results_calculator_n212) );
  BUF_X1 extimating_unit_Results_calculator_U7 ( .A(
        extimating_unit_Results_calculator_n205), .Z(
        extimating_unit_Results_calculator_n209) );
  BUF_X1 extimating_unit_Results_calculator_U6 ( .A(
        extimating_unit_Results_calculator_n205), .Z(
        extimating_unit_Results_calculator_n207) );
  BUF_X1 extimating_unit_Results_calculator_U5 ( .A(
        extimating_unit_Results_calculator_n205), .Z(
        extimating_unit_Results_calculator_n208) );
  BUF_X1 extimating_unit_Results_calculator_U4 ( .A(
        extimating_unit_Results_calculator_n205), .Z(
        extimating_unit_Results_calculator_n210) );
  BUF_X1 extimating_unit_Results_calculator_U3 ( .A(
        extimating_unit_Results_calculator_n205), .Z(
        extimating_unit_Results_calculator_n211) );
  INV_X4 extimating_unit_Results_calculator_U2 ( .A(
        extimating_unit_Results_calculator_n198), .ZN(
        extimating_unit_Results_calculator_n201) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_0__10_ ( .D(
        extimating_unit_Results_calculator_n143), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[10]), .QN(
        extimating_unit_Results_calculator_n77) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_1__10_ ( .D(
        extimating_unit_Results_calculator_n154), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[21]), .QN(
        extimating_unit_Results_calculator_n88) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_1__0_ ( .D(
        extimating_unit_Results_calculator_n144), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[11]), .QN(
        extimating_unit_Results_calculator_n78) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_0__0_ ( .D(
        extimating_unit_Results_calculator_n155), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[0]), .QN(
        extimating_unit_Results_calculator_n89) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_1__0_ ( .D(
        extimating_unit_Results_calculator_n166), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[11]), .QN(
        extimating_unit_Results_calculator_n100) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_0__1_ ( .D(
        extimating_unit_Results_calculator_n156), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[1]), .QN(
        extimating_unit_Results_calculator_n90) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_0__2_ ( .D(
        extimating_unit_Results_calculator_n157), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[2]), .QN(
        extimating_unit_Results_calculator_n91) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_0__4_ ( .D(
        extimating_unit_Results_calculator_n159), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[4]), .QN(
        extimating_unit_Results_calculator_n93) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_0__5_ ( .D(
        extimating_unit_Results_calculator_n160), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[5]), .QN(
        extimating_unit_Results_calculator_n94) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_0__7_ ( .D(
        extimating_unit_Results_calculator_n162), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[7]), .QN(
        extimating_unit_Results_calculator_n96) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_0__8_ ( .D(
        extimating_unit_Results_calculator_n163), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[8]), .QN(
        extimating_unit_Results_calculator_n97) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_0__3_ ( .D(
        extimating_unit_Results_calculator_n158), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[3]), .QN(
        extimating_unit_Results_calculator_n92) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_0__6_ ( .D(
        extimating_unit_Results_calculator_n161), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[6]), .QN(
        extimating_unit_Results_calculator_n95) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_0__9_ ( .D(
        extimating_unit_Results_calculator_n164), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[9]), .QN(
        extimating_unit_Results_calculator_n98) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_0__10_ ( .D(
        extimating_unit_Results_calculator_n165), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[10]), .QN(
        extimating_unit_Results_calculator_n99) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_1__1_ ( .D(
        extimating_unit_Results_calculator_n167), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[12]), .QN(
        extimating_unit_Results_calculator_n101) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_1__2_ ( .D(
        extimating_unit_Results_calculator_n168), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[13]), .QN(
        extimating_unit_Results_calculator_n102) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_1__3_ ( .D(
        extimating_unit_Results_calculator_n169), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[14]), .QN(
        extimating_unit_Results_calculator_n103) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_1__4_ ( .D(
        extimating_unit_Results_calculator_n170), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[15]), .QN(
        extimating_unit_Results_calculator_n104) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_1__5_ ( .D(
        extimating_unit_Results_calculator_n171), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[16]), .QN(
        extimating_unit_Results_calculator_n105) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_1__6_ ( .D(
        extimating_unit_Results_calculator_n172), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[17]), .QN(
        extimating_unit_Results_calculator_n106) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_1__7_ ( .D(
        extimating_unit_Results_calculator_n173), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[18]), .QN(
        extimating_unit_Results_calculator_n107) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_1__8_ ( .D(
        extimating_unit_Results_calculator_n174), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[19]), .QN(
        extimating_unit_Results_calculator_n108) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_1__9_ ( .D(
        extimating_unit_Results_calculator_n175), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[20]), .QN(
        extimating_unit_Results_calculator_n109) );
  DFFR_X1 extimating_unit_Results_calculator_MV0_in_int_reg_1__10_ ( .D(
        extimating_unit_Results_calculator_n176), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV0_out[21]), .QN(
        extimating_unit_Results_calculator_n110) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_1__8_ ( .D(
        extimating_unit_Results_calculator_n152), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[19]), .QN(
        extimating_unit_Results_calculator_n86) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_0__1_ ( .D(
        extimating_unit_Results_calculator_n134), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[1]), .QN(
        extimating_unit_Results_calculator_n68) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_0__4_ ( .D(
        extimating_unit_Results_calculator_n137), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[4]), .QN(
        extimating_unit_Results_calculator_n71) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_0__7_ ( .D(
        extimating_unit_Results_calculator_n140), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[7]), .QN(
        extimating_unit_Results_calculator_n74) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_0__9_ ( .D(
        extimating_unit_Results_calculator_n142), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[9]), .QN(
        extimating_unit_Results_calculator_n76) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_1__1_ ( .D(
        extimating_unit_Results_calculator_n145), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[12]), .QN(
        extimating_unit_Results_calculator_n79) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_1__2_ ( .D(
        extimating_unit_Results_calculator_n146), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[13]), .QN(
        extimating_unit_Results_calculator_n80) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_1__3_ ( .D(
        extimating_unit_Results_calculator_n147), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[14]), .QN(
        extimating_unit_Results_calculator_n81) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_1__4_ ( .D(
        extimating_unit_Results_calculator_n148), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[15]), .QN(
        extimating_unit_Results_calculator_n82) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_1__5_ ( .D(
        extimating_unit_Results_calculator_n149), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[16]), .QN(
        extimating_unit_Results_calculator_n83) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_1__6_ ( .D(
        extimating_unit_Results_calculator_n150), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[17]), .QN(
        extimating_unit_Results_calculator_n84) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_1__7_ ( .D(
        extimating_unit_Results_calculator_n151), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[18]), .QN(
        extimating_unit_Results_calculator_n85) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_1__9_ ( .D(
        extimating_unit_Results_calculator_n153), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[20]), .QN(
        extimating_unit_Results_calculator_n87) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_0__2_ ( .D(
        extimating_unit_Results_calculator_n135), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[2]), .QN(
        extimating_unit_Results_calculator_n69) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_0__3_ ( .D(
        extimating_unit_Results_calculator_n136), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[3]), .QN(
        extimating_unit_Results_calculator_n70) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_0__5_ ( .D(
        extimating_unit_Results_calculator_n138), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[5]), .QN(
        extimating_unit_Results_calculator_n72) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_0__6_ ( .D(
        extimating_unit_Results_calculator_n139), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[6]), .QN(
        extimating_unit_Results_calculator_n73) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_0__8_ ( .D(
        extimating_unit_Results_calculator_n141), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[8]), .QN(
        extimating_unit_Results_calculator_n75) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_1__9_ ( .D(
        extimating_unit_Results_calculator_n197), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[20]), .QN(
        extimating_unit_Results_calculator_n131) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_1__3_ ( .D(
        extimating_unit_Results_calculator_n191), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[14]), .QN(
        extimating_unit_Results_calculator_n125) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_1__5_ ( .D(
        extimating_unit_Results_calculator_n193), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[16]), .QN(
        extimating_unit_Results_calculator_n127) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_1__6_ ( .D(
        extimating_unit_Results_calculator_n194), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[17]), .QN(
        extimating_unit_Results_calculator_n128) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_1__7_ ( .D(
        extimating_unit_Results_calculator_n195), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[18]), .QN(
        extimating_unit_Results_calculator_n129) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_1__8_ ( .D(
        extimating_unit_Results_calculator_n196), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[19]), .QN(
        extimating_unit_Results_calculator_n130) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_1__10_ ( .D(
        extimating_unit_Results_calculator_n199), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[21]), .QN(
        extimating_unit_Results_calculator_n132) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_0__0_ ( .D(
        extimating_unit_Results_calculator_n177), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[0]), .QN(
        extimating_unit_Results_calculator_n111) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_0__1_ ( .D(
        extimating_unit_Results_calculator_n178), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[1]), .QN(
        extimating_unit_Results_calculator_n112) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_0__2_ ( .D(
        extimating_unit_Results_calculator_n179), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[2]), .QN(
        extimating_unit_Results_calculator_n113) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_0__3_ ( .D(
        extimating_unit_Results_calculator_n180), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[3]), .QN(
        extimating_unit_Results_calculator_n114) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_0__4_ ( .D(
        extimating_unit_Results_calculator_n181), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[4]), .QN(
        extimating_unit_Results_calculator_n115) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_0__5_ ( .D(
        extimating_unit_Results_calculator_n182), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[5]), .QN(
        extimating_unit_Results_calculator_n116) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_0__6_ ( .D(
        extimating_unit_Results_calculator_n183), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[6]), .QN(
        extimating_unit_Results_calculator_n117) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_0__7_ ( .D(
        extimating_unit_Results_calculator_n184), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[7]), .QN(
        extimating_unit_Results_calculator_n118) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_0__8_ ( .D(
        extimating_unit_Results_calculator_n185), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[8]), .QN(
        extimating_unit_Results_calculator_n119) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_0__9_ ( .D(
        extimating_unit_Results_calculator_n186), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[9]), .QN(
        extimating_unit_Results_calculator_n120) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_0__10_ ( .D(
        extimating_unit_Results_calculator_n187), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[10]), .QN(
        extimating_unit_Results_calculator_n121) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_1__0_ ( .D(
        extimating_unit_Results_calculator_n188), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[11]), .QN(
        extimating_unit_Results_calculator_n122) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_1__1_ ( .D(
        extimating_unit_Results_calculator_n189), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[12]), .QN(
        extimating_unit_Results_calculator_n123) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_1__2_ ( .D(
        extimating_unit_Results_calculator_n190), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[13]), .QN(
        extimating_unit_Results_calculator_n124) );
  DFFR_X1 extimating_unit_Results_calculator_MV2_in_int_reg_1__4_ ( .D(
        extimating_unit_Results_calculator_n192), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV2_out[15]), .QN(
        extimating_unit_Results_calculator_n126) );
  DFFR_X1 extimating_unit_Results_calculator_MV1_in_int_reg_0__0_ ( .D(
        extimating_unit_Results_calculator_n133), .CK(clk), .RN(
        extimating_unit_Results_calculator_n201), .Q(MV1_out[0]), .QN(
        extimating_unit_Results_calculator_n67) );
  XNOR2_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U12 ( .A(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n10), .B(
        RefPel[0]), .ZN(extimating_unit_Results_calculator_Pel_diff[0]) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U11 ( .A(
        RefPel[0]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n1) );
  NAND2_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U10 ( .A1(
        CurPel[0]), .A2(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n1), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[1]) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U9 ( .A(
        CurPel[1]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n9) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U8 ( .A(
        CurPel[0]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n10) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U7 ( .A(
        CurPel[7]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n3) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U6 ( .A(
        CurPel[6]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n4) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U5 ( .A(
        CurPel[5]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n5) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U4 ( .A(
        CurPel[4]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n6) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U3 ( .A(
        CurPel[3]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n7) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U2 ( .A(
        CurPel[2]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n8) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U1 ( .A(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[8]), .ZN(
        extimating_unit_Results_calculator_Pel_diff[8]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U2_1 ( .A(
        RefPel[1]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n9), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[1]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[2]), .S(
        extimating_unit_Results_calculator_Pel_diff[1]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U2_2 ( .A(
        RefPel[2]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n8), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[2]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[3]), .S(
        extimating_unit_Results_calculator_Pel_diff[2]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U2_3 ( .A(
        RefPel[3]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n7), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[3]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[4]), .S(
        extimating_unit_Results_calculator_Pel_diff[3]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U2_4 ( .A(
        RefPel[4]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n6), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[4]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[5]), .S(
        extimating_unit_Results_calculator_Pel_diff[4]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U2_5 ( .A(
        RefPel[5]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n5), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[5]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[6]), .S(
        extimating_unit_Results_calculator_Pel_diff[5]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U2_6 ( .A(
        RefPel[6]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n4), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[6]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[7]), .S(
        extimating_unit_Results_calculator_Pel_diff[6]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_U2_7 ( .A(
        RefPel[7]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_n3), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[7]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_0_sub_19_carry[8]), .S(
        extimating_unit_Results_calculator_Pel_diff[7]) );
  INV_X1 extimating_unit_Results_calculator_Pel_diff_reg_0_U3 ( .A(
        extimating_unit_Results_calculator_n204), .ZN(
        extimating_unit_Results_calculator_Pel_diff_reg_0_n1) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_0_Q_int_reg_7_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[7]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[7]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_0_Q_int_reg_8_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[8]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[8]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_0_Q_int_reg_6_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[6]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[6]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_0_Q_int_reg_5_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[5]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[5]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_0_Q_int_reg_4_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[4]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[4]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_0_Q_int_reg_3_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[3]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[3]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_0_Q_int_reg_2_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[2]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[2]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_0_Q_int_reg_1_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[1]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[1]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_0_Q_int_reg_0_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[0]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[0]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_0_U39 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[7]), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_0_n7), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[8]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n14) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U38 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n14), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[7]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_0_U37 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[6]), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_0_n6), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[8]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n15) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U36 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n15), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[6]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_0_U35 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[5]), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_0_n5), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[8]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n16) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U34 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n16), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[5]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_0_U33 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[4]), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_0_n4), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[8]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n17) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U32 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n17), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[4]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_0_U31 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[3]), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_0_n3), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[8]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n18) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U30 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n18), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[3]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_0_U29 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[2]), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_0_n2), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[8]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n19) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U28 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n19), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[2]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_0_U27 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[1]), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_0_n1), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[8]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n20) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U26 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n20), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[1]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_0_U25 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[0]), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n38), .B1(
        extimating_unit_Results_calculator_Pel_diff_samp[0]), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[8]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n21) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U24 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n21), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[0]) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U23 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[7]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n29) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U22 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[6]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n28) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U21 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[5]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n27) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U20 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[4]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n26) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U19 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[3]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n25) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U18 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[2]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n24) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U17 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[1]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n23) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U16 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[0]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n22) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_0_U15 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[8]), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n38) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_0_U14 ( .A1(
        extimating_unit_Results_calculator_Abs_X_0_n28), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n12), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n13) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_0_U13 ( .A1(
        extimating_unit_Results_calculator_Abs_X_0_n27), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n11), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n12) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_0_U12 ( .A1(
        extimating_unit_Results_calculator_Abs_X_0_n26), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n10), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n11) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_0_U11 ( .A1(
        extimating_unit_Results_calculator_Abs_X_0_n25), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n9), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n10) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_0_U10 ( .A1(
        extimating_unit_Results_calculator_Abs_X_0_n24), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n8), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n9) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_0_U9 ( .A1(
        extimating_unit_Results_calculator_Abs_X_0_n23), .A2(
        extimating_unit_Results_calculator_Abs_X_0_n22), .ZN(
        extimating_unit_Results_calculator_Abs_X_0_n8) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_0_U8 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n29), .B(
        extimating_unit_Results_calculator_Abs_X_0_n13), .Z(
        extimating_unit_Results_calculator_Abs_X_0_n7) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_0_U7 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n28), .B(
        extimating_unit_Results_calculator_Abs_X_0_n12), .Z(
        extimating_unit_Results_calculator_Abs_X_0_n6) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_0_U6 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n27), .B(
        extimating_unit_Results_calculator_Abs_X_0_n11), .Z(
        extimating_unit_Results_calculator_Abs_X_0_n5) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_0_U5 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n26), .B(
        extimating_unit_Results_calculator_Abs_X_0_n10), .Z(
        extimating_unit_Results_calculator_Abs_X_0_n4) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_0_U4 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n25), .B(
        extimating_unit_Results_calculator_Abs_X_0_n9), .Z(
        extimating_unit_Results_calculator_Abs_X_0_n3) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_0_U3 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n24), .B(
        extimating_unit_Results_calculator_Abs_X_0_n8), .Z(
        extimating_unit_Results_calculator_Abs_X_0_n2) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_0_U2 ( .A(
        extimating_unit_Results_calculator_Abs_X_0_n23), .B(
        extimating_unit_Results_calculator_Abs_X_0_n22), .Z(
        extimating_unit_Results_calculator_Abs_X_0_n1) );
  INV_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_U3 ( .A(
        extimating_unit_Results_calculator_n202), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_n1) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_Q_int_reg_7_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[7]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[7]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_Q_int_reg_6_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[6]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[6]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_Q_int_reg_5_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[5]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[5]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_Q_int_reg_4_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[4]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[4]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_Q_int_reg_3_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[3]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[3]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_Q_int_reg_2_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[2]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[2]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_Q_int_reg_0_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[0]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[0]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_Q_int_reg_1_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[1]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_0_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[1]) );
  XNOR2_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U12 ( .A(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n10), .B(
        RefPel[8]), .ZN(extimating_unit_Results_calculator_Pel_diff[9]) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U11 ( .A(
        RefPel[8]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n1) );
  NAND2_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U10 ( .A1(
        CurPel[8]), .A2(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n1), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[1]) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U9 ( .A(
        CurPel[9]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n9) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U8 ( .A(
        CurPel[8]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n10) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U7 ( .A(
        CurPel[15]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n3) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U6 ( .A(
        CurPel[14]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n4) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U5 ( .A(
        CurPel[13]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n5) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U4 ( .A(
        CurPel[12]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n6) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U3 ( .A(
        CurPel[11]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n7) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U2 ( .A(
        CurPel[10]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n8) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U1 ( .A(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[8]), .ZN(
        extimating_unit_Results_calculator_Pel_diff[17]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U2_1 ( .A(
        RefPel[9]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n9), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[1]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[2]), .S(
        extimating_unit_Results_calculator_Pel_diff[10]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U2_2 ( .A(
        RefPel[10]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n8), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[2]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[3]), .S(
        extimating_unit_Results_calculator_Pel_diff[11]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U2_3 ( .A(
        RefPel[11]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n7), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[3]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[4]), .S(
        extimating_unit_Results_calculator_Pel_diff[12]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U2_4 ( .A(
        RefPel[12]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n6), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[4]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[5]), .S(
        extimating_unit_Results_calculator_Pel_diff[13]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U2_5 ( .A(
        RefPel[13]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n5), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[5]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[6]), .S(
        extimating_unit_Results_calculator_Pel_diff[14]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U2_6 ( .A(
        RefPel[14]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n4), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[6]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[7]), .S(
        extimating_unit_Results_calculator_Pel_diff[15]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_U2_7 ( .A(
        RefPel[15]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_n3), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[7]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_1_sub_19_carry[8]), .S(
        extimating_unit_Results_calculator_Pel_diff[16]) );
  INV_X1 extimating_unit_Results_calculator_Pel_diff_reg_1_U3 ( .A(
        extimating_unit_Results_calculator_n204), .ZN(
        extimating_unit_Results_calculator_Pel_diff_reg_1_n1) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_1_Q_int_reg_0_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[9]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[9]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_1_Q_int_reg_1_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[10]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[10]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_1_Q_int_reg_2_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[11]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[11]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_1_Q_int_reg_3_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[12]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[12]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_1_Q_int_reg_4_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[13]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[13]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_1_Q_int_reg_5_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[14]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[14]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_1_Q_int_reg_6_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[15]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[15]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_1_Q_int_reg_7_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[16]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[16]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_1_Q_int_reg_8_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[17]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[17]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_1_U39 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[16]), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_1_n7), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[17]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n46) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U38 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n46), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[15]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_1_U37 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[15]), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_1_n6), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[17]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n45) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U36 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n45), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[14]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_1_U35 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[14]), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_1_n5), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[17]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n44) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U34 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n44), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[13]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_1_U33 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[13]), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_1_n4), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[17]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n43) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U32 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n43), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[12]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_1_U31 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[12]), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_1_n3), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[17]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n42) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U30 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n42), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[11]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_1_U29 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[11]), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_1_n2), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[17]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n41) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U28 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n41), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[10]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_1_U27 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[10]), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_1_n1), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[17]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n40) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U26 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n40), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[9]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_1_U25 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[9]), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n38), .B1(
        extimating_unit_Results_calculator_Pel_diff_samp[9]), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[17]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n39) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U24 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n39), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[8]) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U23 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[16]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n29) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U22 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[15]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n28) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U21 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[14]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n27) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U20 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[13]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n26) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U19 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[12]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n25) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U18 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[11]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n24) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U17 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[10]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n23) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U16 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[9]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n22) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_1_U15 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[17]), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n38) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_1_U14 ( .A1(
        extimating_unit_Results_calculator_Abs_X_1_n28), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n12), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n13) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_1_U13 ( .A1(
        extimating_unit_Results_calculator_Abs_X_1_n27), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n11), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n12) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_1_U12 ( .A1(
        extimating_unit_Results_calculator_Abs_X_1_n26), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n10), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n11) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_1_U11 ( .A1(
        extimating_unit_Results_calculator_Abs_X_1_n25), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n9), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n10) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_1_U10 ( .A1(
        extimating_unit_Results_calculator_Abs_X_1_n24), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n8), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n9) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_1_U9 ( .A1(
        extimating_unit_Results_calculator_Abs_X_1_n23), .A2(
        extimating_unit_Results_calculator_Abs_X_1_n22), .ZN(
        extimating_unit_Results_calculator_Abs_X_1_n8) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_1_U8 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n29), .B(
        extimating_unit_Results_calculator_Abs_X_1_n13), .Z(
        extimating_unit_Results_calculator_Abs_X_1_n7) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_1_U7 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n28), .B(
        extimating_unit_Results_calculator_Abs_X_1_n12), .Z(
        extimating_unit_Results_calculator_Abs_X_1_n6) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_1_U6 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n27), .B(
        extimating_unit_Results_calculator_Abs_X_1_n11), .Z(
        extimating_unit_Results_calculator_Abs_X_1_n5) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_1_U5 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n26), .B(
        extimating_unit_Results_calculator_Abs_X_1_n10), .Z(
        extimating_unit_Results_calculator_Abs_X_1_n4) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_1_U4 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n25), .B(
        extimating_unit_Results_calculator_Abs_X_1_n9), .Z(
        extimating_unit_Results_calculator_Abs_X_1_n3) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_1_U3 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n24), .B(
        extimating_unit_Results_calculator_Abs_X_1_n8), .Z(
        extimating_unit_Results_calculator_Abs_X_1_n2) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_1_U2 ( .A(
        extimating_unit_Results_calculator_Abs_X_1_n23), .B(
        extimating_unit_Results_calculator_Abs_X_1_n22), .Z(
        extimating_unit_Results_calculator_Abs_X_1_n1) );
  INV_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_U3 ( .A(
        extimating_unit_Results_calculator_n204), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_n1) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_Q_int_reg_0_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[8]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[8]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_Q_int_reg_1_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[9]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[9]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_Q_int_reg_2_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[10]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[10]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_Q_int_reg_3_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[11]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[11]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_Q_int_reg_4_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[12]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[12]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_Q_int_reg_5_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[13]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[13]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_Q_int_reg_6_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[14]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[14]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_Q_int_reg_7_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[15]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_1_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[15]) );
  XNOR2_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U12 ( .A(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n10), .B(
        RefPel[16]), .ZN(extimating_unit_Results_calculator_Pel_diff[18]) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U11 ( .A(
        RefPel[16]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n1) );
  NAND2_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U10 ( .A1(
        CurPel[16]), .A2(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n1), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[1]) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U9 ( .A(
        CurPel[17]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n9) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U8 ( .A(
        CurPel[16]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n10) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U7 ( .A(
        CurPel[23]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n3) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U6 ( .A(
        CurPel[22]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n4) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U5 ( .A(
        CurPel[21]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n5) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U4 ( .A(
        CurPel[20]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n6) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U3 ( .A(
        CurPel[19]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n7) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U2 ( .A(
        CurPel[18]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n8) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U1 ( .A(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[8]), .ZN(
        extimating_unit_Results_calculator_Pel_diff[26]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U2_1 ( .A(
        RefPel[17]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n9), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[1]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[2]), .S(
        extimating_unit_Results_calculator_Pel_diff[19]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U2_2 ( .A(
        RefPel[18]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n8), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[2]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[3]), .S(
        extimating_unit_Results_calculator_Pel_diff[20]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U2_3 ( .A(
        RefPel[19]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n7), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[3]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[4]), .S(
        extimating_unit_Results_calculator_Pel_diff[21]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U2_4 ( .A(
        RefPel[20]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n6), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[4]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[5]), .S(
        extimating_unit_Results_calculator_Pel_diff[22]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U2_5 ( .A(
        RefPel[21]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n5), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[5]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[6]), .S(
        extimating_unit_Results_calculator_Pel_diff[23]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U2_6 ( .A(
        RefPel[22]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n4), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[6]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[7]), .S(
        extimating_unit_Results_calculator_Pel_diff[24]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_U2_7 ( .A(
        RefPel[23]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_n3), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[7]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_2_sub_19_carry[8]), .S(
        extimating_unit_Results_calculator_Pel_diff[25]) );
  INV_X1 extimating_unit_Results_calculator_Pel_diff_reg_2_U3 ( .A(
        extimating_unit_Results_calculator_n204), .ZN(
        extimating_unit_Results_calculator_Pel_diff_reg_2_n1) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_2_Q_int_reg_0_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[18]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[18]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_2_Q_int_reg_1_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[19]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[19]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_2_Q_int_reg_2_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[20]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[20]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_2_Q_int_reg_3_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[21]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[21]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_2_Q_int_reg_4_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[22]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[22]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_2_Q_int_reg_5_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[23]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[23]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_2_Q_int_reg_6_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[24]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[24]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_2_Q_int_reg_7_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[25]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[25]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_2_Q_int_reg_8_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[26]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[26]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_2_U39 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[25]), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_2_n7), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[26]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n46) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U38 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n46), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[23]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_2_U37 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[24]), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_2_n6), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[26]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n45) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U36 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n45), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[22]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_2_U35 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[23]), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_2_n5), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[26]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n44) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U34 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n44), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[21]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_2_U33 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[22]), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_2_n4), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[26]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n43) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U32 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n43), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[20]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_2_U31 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[21]), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_2_n3), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[26]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n42) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U30 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n42), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[19]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_2_U29 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[20]), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_2_n2), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[26]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n41) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U28 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n41), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[18]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_2_U27 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[19]), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_2_n1), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[26]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n40) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U26 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n40), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[17]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_2_U25 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[18]), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n38), .B1(
        extimating_unit_Results_calculator_Pel_diff_samp[18]), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[26]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n39) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U24 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n39), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[16]) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U23 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[25]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n29) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U22 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[24]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n28) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U21 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[23]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n27) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U20 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[22]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n26) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U19 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[21]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n25) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U18 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[20]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n24) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U17 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[19]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n23) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U16 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[18]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n22) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_2_U15 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[26]), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n38) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_2_U14 ( .A1(
        extimating_unit_Results_calculator_Abs_X_2_n28), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n12), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n13) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_2_U13 ( .A1(
        extimating_unit_Results_calculator_Abs_X_2_n27), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n11), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n12) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_2_U12 ( .A1(
        extimating_unit_Results_calculator_Abs_X_2_n26), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n10), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n11) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_2_U11 ( .A1(
        extimating_unit_Results_calculator_Abs_X_2_n25), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n9), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n10) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_2_U10 ( .A1(
        extimating_unit_Results_calculator_Abs_X_2_n24), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n8), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n9) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_2_U9 ( .A1(
        extimating_unit_Results_calculator_Abs_X_2_n23), .A2(
        extimating_unit_Results_calculator_Abs_X_2_n22), .ZN(
        extimating_unit_Results_calculator_Abs_X_2_n8) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_2_U8 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n29), .B(
        extimating_unit_Results_calculator_Abs_X_2_n13), .Z(
        extimating_unit_Results_calculator_Abs_X_2_n7) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_2_U7 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n28), .B(
        extimating_unit_Results_calculator_Abs_X_2_n12), .Z(
        extimating_unit_Results_calculator_Abs_X_2_n6) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_2_U6 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n27), .B(
        extimating_unit_Results_calculator_Abs_X_2_n11), .Z(
        extimating_unit_Results_calculator_Abs_X_2_n5) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_2_U5 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n26), .B(
        extimating_unit_Results_calculator_Abs_X_2_n10), .Z(
        extimating_unit_Results_calculator_Abs_X_2_n4) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_2_U4 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n25), .B(
        extimating_unit_Results_calculator_Abs_X_2_n9), .Z(
        extimating_unit_Results_calculator_Abs_X_2_n3) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_2_U3 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n24), .B(
        extimating_unit_Results_calculator_Abs_X_2_n8), .Z(
        extimating_unit_Results_calculator_Abs_X_2_n2) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_2_U2 ( .A(
        extimating_unit_Results_calculator_Abs_X_2_n23), .B(
        extimating_unit_Results_calculator_Abs_X_2_n22), .Z(
        extimating_unit_Results_calculator_Abs_X_2_n1) );
  INV_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_U3 ( .A(
        extimating_unit_Results_calculator_n204), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_n1) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_Q_int_reg_0_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[16]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[16]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_Q_int_reg_1_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[17]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[17]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_Q_int_reg_2_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[18]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[18]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_Q_int_reg_3_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[19]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[19]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_Q_int_reg_4_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[20]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[20]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_Q_int_reg_5_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[21]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[21]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_Q_int_reg_6_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[22]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[22]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_Q_int_reg_7_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[23]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_2_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[23]) );
  XNOR2_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U12 ( .A(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n10), .B(
        RefPel[24]), .ZN(extimating_unit_Results_calculator_Pel_diff[27]) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U11 ( .A(
        RefPel[24]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n1) );
  NAND2_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U10 ( .A1(
        CurPel[24]), .A2(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n1), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[1]) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U9 ( .A(
        CurPel[25]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n9) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U8 ( .A(
        CurPel[24]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n10) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U7 ( .A(
        CurPel[31]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n3) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U6 ( .A(
        CurPel[30]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n4) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U5 ( .A(
        CurPel[29]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n5) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U4 ( .A(
        CurPel[28]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n6) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U3 ( .A(
        CurPel[27]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n7) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U2 ( .A(
        CurPel[26]), .ZN(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n8) );
  INV_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U1 ( .A(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[8]), .ZN(
        extimating_unit_Results_calculator_Pel_diff[35]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U2_1 ( .A(
        RefPel[25]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n9), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[1]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[2]), .S(
        extimating_unit_Results_calculator_Pel_diff[28]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U2_2 ( .A(
        RefPel[26]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n8), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[2]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[3]), .S(
        extimating_unit_Results_calculator_Pel_diff[29]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U2_3 ( .A(
        RefPel[27]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n7), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[3]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[4]), .S(
        extimating_unit_Results_calculator_Pel_diff[30]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U2_4 ( .A(
        RefPel[28]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n6), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[4]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[5]), .S(
        extimating_unit_Results_calculator_Pel_diff[31]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U2_5 ( .A(
        RefPel[29]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n5), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[5]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[6]), .S(
        extimating_unit_Results_calculator_Pel_diff[32]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U2_6 ( .A(
        RefPel[30]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n4), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[6]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[7]), .S(
        extimating_unit_Results_calculator_Pel_diff[33]) );
  FA_X1 extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_U2_7 ( .A(
        RefPel[31]), .B(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_n3), .CI(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[7]), .CO(
        extimating_unit_Results_calculator_Pel_sub_X_3_sub_19_carry[8]), .S(
        extimating_unit_Results_calculator_Pel_diff[34]) );
  INV_X1 extimating_unit_Results_calculator_Pel_diff_reg_3_U3 ( .A(
        extimating_unit_Results_calculator_n203), .ZN(
        extimating_unit_Results_calculator_Pel_diff_reg_3_n1) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_3_Q_int_reg_0_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[27]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[27]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_3_Q_int_reg_1_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[28]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[28]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_3_Q_int_reg_2_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[29]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[29]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_3_Q_int_reg_3_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[30]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[30]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_3_Q_int_reg_4_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[31]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[31]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_3_Q_int_reg_5_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[32]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[32]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_3_Q_int_reg_6_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[33]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[33]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_3_Q_int_reg_7_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[34]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[34]) );
  DFFR_X1 extimating_unit_Results_calculator_Pel_diff_reg_3_Q_int_reg_8_ ( .D(
        extimating_unit_Results_calculator_Pel_diff[35]), .CK(clk), .RN(
        extimating_unit_Results_calculator_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_Pel_diff_samp[35]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_3_U39 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[34]), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_3_n7), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[35]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n46) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U38 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n46), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[31]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_3_U37 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[33]), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_3_n6), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[35]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n45) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U36 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n45), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[30]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_3_U35 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[32]), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_3_n5), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[35]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n44) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U34 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n44), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[29]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_3_U33 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[31]), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_3_n4), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[35]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n43) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U32 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n43), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[28]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_3_U31 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[30]), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_3_n3), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[35]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n42) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U30 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n42), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[27]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_3_U29 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[29]), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_3_n2), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[35]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n41) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U28 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n41), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[26]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_3_U27 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[28]), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n38), .B1(
        extimating_unit_Results_calculator_Abs_X_3_n1), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[35]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n40) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U26 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n40), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[25]) );
  AOI22_X1 extimating_unit_Results_calculator_Abs_X_3_U25 ( .A1(
        extimating_unit_Results_calculator_Pel_diff_samp[27]), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n38), .B1(
        extimating_unit_Results_calculator_Pel_diff_samp[27]), .B2(
        extimating_unit_Results_calculator_Pel_diff_samp[35]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n39) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U24 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n39), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff[24]) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U23 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[34]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n29) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U22 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[33]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n28) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U21 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[32]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n27) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U20 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[31]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n26) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U19 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[30]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n25) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U18 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[29]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n24) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U17 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[28]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n23) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U16 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[27]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n22) );
  INV_X1 extimating_unit_Results_calculator_Abs_X_3_U15 ( .A(
        extimating_unit_Results_calculator_Pel_diff_samp[35]), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n38) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_3_U14 ( .A1(
        extimating_unit_Results_calculator_Abs_X_3_n28), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n12), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n13) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_3_U13 ( .A1(
        extimating_unit_Results_calculator_Abs_X_3_n27), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n11), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n12) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_3_U12 ( .A1(
        extimating_unit_Results_calculator_Abs_X_3_n26), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n10), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n11) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_3_U11 ( .A1(
        extimating_unit_Results_calculator_Abs_X_3_n25), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n9), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n10) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_3_U10 ( .A1(
        extimating_unit_Results_calculator_Abs_X_3_n24), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n8), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n9) );
  AND2_X1 extimating_unit_Results_calculator_Abs_X_3_U9 ( .A1(
        extimating_unit_Results_calculator_Abs_X_3_n23), .A2(
        extimating_unit_Results_calculator_Abs_X_3_n22), .ZN(
        extimating_unit_Results_calculator_Abs_X_3_n8) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_3_U8 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n29), .B(
        extimating_unit_Results_calculator_Abs_X_3_n13), .Z(
        extimating_unit_Results_calculator_Abs_X_3_n7) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_3_U7 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n28), .B(
        extimating_unit_Results_calculator_Abs_X_3_n12), .Z(
        extimating_unit_Results_calculator_Abs_X_3_n6) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_3_U6 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n27), .B(
        extimating_unit_Results_calculator_Abs_X_3_n11), .Z(
        extimating_unit_Results_calculator_Abs_X_3_n5) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_3_U5 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n26), .B(
        extimating_unit_Results_calculator_Abs_X_3_n10), .Z(
        extimating_unit_Results_calculator_Abs_X_3_n4) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_3_U4 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n25), .B(
        extimating_unit_Results_calculator_Abs_X_3_n9), .Z(
        extimating_unit_Results_calculator_Abs_X_3_n3) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_3_U3 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n24), .B(
        extimating_unit_Results_calculator_Abs_X_3_n8), .Z(
        extimating_unit_Results_calculator_Abs_X_3_n2) );
  XOR2_X1 extimating_unit_Results_calculator_Abs_X_3_U2 ( .A(
        extimating_unit_Results_calculator_Abs_X_3_n23), .B(
        extimating_unit_Results_calculator_Abs_X_3_n22), .Z(
        extimating_unit_Results_calculator_Abs_X_3_n1) );
  INV_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_U3 ( .A(
        extimating_unit_Results_calculator_n204), .ZN(
        extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_n1) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_Q_int_reg_0_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[24]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[24]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_Q_int_reg_1_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[25]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[25]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_Q_int_reg_2_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[26]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[26]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_Q_int_reg_3_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[27]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[27]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_Q_int_reg_4_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[28]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[28]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_Q_int_reg_5_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[29]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[29]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_Q_int_reg_6_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[30]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[30]) );
  DFFR_X1 extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_Q_int_reg_7_ ( 
        .D(extimating_unit_Results_calculator_Abs_Pel_diff[31]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Abs_Pel_diff_reg_3_n1), .Q(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[31]) );
  XOR2_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_U2 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[8]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[0]), .Z(
        extimating_unit_Results_calculator_PelAdd_stage1_out[0]) );
  AND2_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_U1 ( 
        .A1(extimating_unit_Results_calculator_ABs_Pel_diff_samp[8]), .A2(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[0]), .ZN(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_n1) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_U1_1 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[1]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[9]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_n1), .CO(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_carry[2]), 
        .S(extimating_unit_Results_calculator_PelAdd_stage1_out[1]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_U1_2 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[2]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[10]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_carry[2]), 
        .CO(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_carry[3]), 
        .S(extimating_unit_Results_calculator_PelAdd_stage1_out[2]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_U1_3 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[3]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[11]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_carry[3]), 
        .CO(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_carry[4]), 
        .S(extimating_unit_Results_calculator_PelAdd_stage1_out[3]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_U1_4 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[4]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[12]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_carry[4]), 
        .CO(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_carry[5]), 
        .S(extimating_unit_Results_calculator_PelAdd_stage1_out[4]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_U1_5 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[5]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[13]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_carry[5]), 
        .CO(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_carry[6]), 
        .S(extimating_unit_Results_calculator_PelAdd_stage1_out[5]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_U1_6 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[6]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[14]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_carry[6]), 
        .CO(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_carry[7]), 
        .S(extimating_unit_Results_calculator_PelAdd_stage1_out[6]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_U1_7 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[7]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[15]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_0_add_23_carry[7]), 
        .CO(extimating_unit_Results_calculator_PelAdd_stage1_out[8]), .S(
        extimating_unit_Results_calculator_PelAdd_stage1_out[7]) );
  INV_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_U3 ( .A(
        extimating_unit_Results_calculator_n203), .ZN(
        extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_n1) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_Q_int_reg_0_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[0]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[0]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_Q_int_reg_1_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[1]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[1]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_Q_int_reg_2_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[2]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[2]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_Q_int_reg_3_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[3]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[3]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_Q_int_reg_4_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[4]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[4]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_Q_int_reg_5_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[5]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[5]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_Q_int_reg_6_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[6]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[6]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_Q_int_reg_7_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[7]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[7]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_Q_int_reg_8_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[8]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_0_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[8]) );
  XOR2_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_U2 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[24]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[16]), .Z(
        extimating_unit_Results_calculator_PelAdd_stage1_out[9]) );
  AND2_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_U1 ( 
        .A1(extimating_unit_Results_calculator_ABs_Pel_diff_samp[24]), .A2(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[16]), .ZN(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_n1) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_U1_1 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[17]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[25]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_n1), .CO(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_carry[2]), 
        .S(extimating_unit_Results_calculator_PelAdd_stage1_out[10]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_U1_2 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[18]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[26]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_carry[2]), 
        .CO(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_carry[3]), 
        .S(extimating_unit_Results_calculator_PelAdd_stage1_out[11]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_U1_3 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[19]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[27]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_carry[3]), 
        .CO(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_carry[4]), 
        .S(extimating_unit_Results_calculator_PelAdd_stage1_out[12]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_U1_4 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[20]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[28]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_carry[4]), 
        .CO(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_carry[5]), 
        .S(extimating_unit_Results_calculator_PelAdd_stage1_out[13]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_U1_5 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[21]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[29]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_carry[5]), 
        .CO(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_carry[6]), 
        .S(extimating_unit_Results_calculator_PelAdd_stage1_out[14]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_U1_6 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[22]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[30]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_carry[6]), 
        .CO(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_carry[7]), 
        .S(extimating_unit_Results_calculator_PelAdd_stage1_out[15]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_U1_7 ( .A(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[23]), .B(
        extimating_unit_Results_calculator_ABs_Pel_diff_samp[31]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage1_X_1_add_23_carry[7]), 
        .CO(extimating_unit_Results_calculator_PelAdd_stage1_out[17]), .S(
        extimating_unit_Results_calculator_PelAdd_stage1_out[16]) );
  INV_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_U3 ( .A(
        extimating_unit_Results_calculator_n203), .ZN(
        extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_n1) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_Q_int_reg_0_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[9]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[9]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_Q_int_reg_1_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[10]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[10]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_Q_int_reg_2_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[11]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[11]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_Q_int_reg_3_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[12]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[12]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_Q_int_reg_4_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[13]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[13]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_Q_int_reg_5_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[14]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[14]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_Q_int_reg_6_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[15]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[15]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_Q_int_reg_7_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[16]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[16]) );
  DFFR_X1 extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_Q_int_reg_8_ ( 
        .D(extimating_unit_Results_calculator_PelAdd_stage1_out[17]), .CK(clk), 
        .RN(extimating_unit_Results_calculator_PelAdd_stage1_out_reg_1_n1), 
        .Q(extimating_unit_Results_calculator_PelAdd_stage1_out_samp[17]) );
  XOR2_X1 extimating_unit_Results_calculator_PelAdd_stage2_add_23_U2 ( .A(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[9]), .B(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[0]), .Z(
        extimating_unit_Results_calculator_PelAdd_out[0]) );
  AND2_X1 extimating_unit_Results_calculator_PelAdd_stage2_add_23_U1 ( .A1(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[9]), .A2(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[0]), .ZN(
        extimating_unit_Results_calculator_PelAdd_stage2_add_23_n1) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage2_add_23_U1_1 ( .A(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[1]), .B(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[10]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage2_add_23_n1), .CO(
        extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[2]), .S(
        extimating_unit_Results_calculator_PelAdd_out[1]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage2_add_23_U1_2 ( .A(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[2]), .B(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[11]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[2]), 
        .CO(extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[3]), 
        .S(extimating_unit_Results_calculator_PelAdd_out[2]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage2_add_23_U1_3 ( .A(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[3]), .B(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[12]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[3]), 
        .CO(extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[4]), 
        .S(extimating_unit_Results_calculator_PelAdd_out[3]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage2_add_23_U1_4 ( .A(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[4]), .B(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[13]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[4]), 
        .CO(extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[5]), 
        .S(extimating_unit_Results_calculator_PelAdd_out[4]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage2_add_23_U1_5 ( .A(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[5]), .B(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[14]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[5]), 
        .CO(extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[6]), 
        .S(extimating_unit_Results_calculator_PelAdd_out[5]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage2_add_23_U1_6 ( .A(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[6]), .B(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[15]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[6]), 
        .CO(extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[7]), 
        .S(extimating_unit_Results_calculator_PelAdd_out[6]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage2_add_23_U1_7 ( .A(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[7]), .B(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[16]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[7]), 
        .CO(extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[8]), 
        .S(extimating_unit_Results_calculator_PelAdd_out[7]) );
  FA_X1 extimating_unit_Results_calculator_PelAdd_stage2_add_23_U1_8 ( .A(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[8]), .B(
        extimating_unit_Results_calculator_PelAdd_stage1_out_samp[17]), .CI(
        extimating_unit_Results_calculator_PelAdd_stage2_add_23_carry[8]), 
        .CO(extimating_unit_Results_calculator_PelAdd_out[9]), .S(
        extimating_unit_Results_calculator_PelAdd_out[8]) );
  INV_X1 extimating_unit_Results_calculator_CurRowSAD_reg_U3 ( .A(
        extimating_unit_Results_calculator_n202), .ZN(
        extimating_unit_Results_calculator_CurRowSAD_reg_n1) );
  DFFR_X1 extimating_unit_Results_calculator_CurRowSAD_reg_Q_int_reg_8_ ( .D(
        extimating_unit_Results_calculator_PelAdd_out[8]), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurRowSAD_reg_n1), .Q(
        extimating_unit_Results_calculator_CurRowSAD[8]) );
  DFFR_X1 extimating_unit_Results_calculator_CurRowSAD_reg_Q_int_reg_9_ ( .D(
        extimating_unit_Results_calculator_PelAdd_out[9]), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurRowSAD_reg_n1), .Q(
        extimating_unit_Results_calculator_CurRowSAD[9]) );
  DFFR_X1 extimating_unit_Results_calculator_CurRowSAD_reg_Q_int_reg_7_ ( .D(
        extimating_unit_Results_calculator_PelAdd_out[7]), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurRowSAD_reg_n1), .Q(
        extimating_unit_Results_calculator_CurRowSAD[7]) );
  DFFR_X1 extimating_unit_Results_calculator_CurRowSAD_reg_Q_int_reg_6_ ( .D(
        extimating_unit_Results_calculator_PelAdd_out[6]), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurRowSAD_reg_n1), .Q(
        extimating_unit_Results_calculator_CurRowSAD[6]) );
  DFFR_X1 extimating_unit_Results_calculator_CurRowSAD_reg_Q_int_reg_5_ ( .D(
        extimating_unit_Results_calculator_PelAdd_out[5]), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurRowSAD_reg_n1), .Q(
        extimating_unit_Results_calculator_CurRowSAD[5]) );
  DFFR_X1 extimating_unit_Results_calculator_CurRowSAD_reg_Q_int_reg_4_ ( .D(
        extimating_unit_Results_calculator_PelAdd_out[4]), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurRowSAD_reg_n1), .Q(
        extimating_unit_Results_calculator_CurRowSAD[4]) );
  DFFR_X1 extimating_unit_Results_calculator_CurRowSAD_reg_Q_int_reg_3_ ( .D(
        extimating_unit_Results_calculator_PelAdd_out[3]), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurRowSAD_reg_n1), .Q(
        extimating_unit_Results_calculator_CurRowSAD[3]) );
  DFFR_X1 extimating_unit_Results_calculator_CurRowSAD_reg_Q_int_reg_2_ ( .D(
        extimating_unit_Results_calculator_PelAdd_out[2]), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurRowSAD_reg_n1), .Q(
        extimating_unit_Results_calculator_CurRowSAD[2]) );
  DFFR_X1 extimating_unit_Results_calculator_CurRowSAD_reg_Q_int_reg_1_ ( .D(
        extimating_unit_Results_calculator_PelAdd_out[1]), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurRowSAD_reg_n1), .Q(
        extimating_unit_Results_calculator_CurRowSAD[1]) );
  DFFR_X1 extimating_unit_Results_calculator_CurRowSAD_reg_Q_int_reg_0_ ( .D(
        extimating_unit_Results_calculator_PelAdd_out[0]), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurRowSAD_reg_n1), .Q(
        extimating_unit_Results_calculator_CurRowSAD[0]) );
  INV_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U21 ( .A(SAD_tmp_RST), 
        .ZN(extimating_unit_Results_calculator_SAD_tmp_reg_n19) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U20 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_0_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n18) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U19 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_1_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n17) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U18 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_2_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n16) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U17 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_3_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n15) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U16 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_4_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n14) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U15 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_5_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n13) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U14 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_6_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n12) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U13 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_7_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n11) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U12 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_8_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n10) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U11 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_9_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n9) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U10 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_10_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n8) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U9 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_11_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n7) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U8 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_12_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n6) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U7 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_13_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n5) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U6 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_14_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n4) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U5 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_15_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n3) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U4 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_16_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n2) );
  AND2_X1 extimating_unit_Results_calculator_SAD_tmp_reg_U3 ( .A1(
        extimating_unit_Results_calculator_CurSAD_tmp_17_), .A2(
        extimating_unit_Results_calculator_SAD_tmp_reg_n19), .ZN(
        extimating_unit_Results_calculator_SAD_tmp_reg_n1) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_17_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n1), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[17]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_16_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n2), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[16]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_15_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n3), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[15]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_14_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n4), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[14]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_13_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n5), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[13]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_12_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n6), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[12]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_11_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n7), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[11]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_10_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n8), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[10]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_9_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n9), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[9]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_8_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n10), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[8]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_7_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n11), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[7]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_6_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n12), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[6]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_5_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n13), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[5]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_4_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n14), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[4]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_3_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n15), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[3]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_2_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n16), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[2]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_1_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n17), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[1]) );
  DFF_X1 extimating_unit_Results_calculator_SAD_tmp_reg_Q_int_reg_0_ ( .D(
        extimating_unit_Results_calculator_SAD_tmp_reg_n18), .CK(clk), .Q(
        extimating_unit_Results_calculator_SAD_tmp[0]) );
  INV_X1 extimating_unit_Results_calculator_CurSAD_reg_U3 ( .A(
        extimating_unit_Results_calculator_n202), .ZN(
        extimating_unit_Results_calculator_CurSAD_reg_n1) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_17_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_17_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[17]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_16_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_16_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[16]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_15_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_15_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[15]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_14_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_14_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[14]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_13_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_13_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[13]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_12_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_12_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[12]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_11_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_11_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[11]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_10_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_10_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[10]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_9_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_9_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[9]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_8_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_8_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[8]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_7_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_7_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[7]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_6_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_6_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[6]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_5_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_5_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[5]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_4_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_4_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[4]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_3_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_3_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[3]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_2_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_2_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[2]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_1_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_1_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[1]) );
  DFFR_X1 extimating_unit_Results_calculator_CurSAD_reg_Q_int_reg_0_ ( .D(
        extimating_unit_Results_calculator_CurSAD_tmp_0_), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurSAD_reg_n1), .Q(CurSAD[0]) );
  OAI22_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U157 ( 
        .A1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n134), 
        .A2(CurSAD[16]), .B1(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n133), .B2(
        CurSAD[17]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n197) );
  AND2_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U156 ( 
        .A1(CurSAD[17]), .A2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n133), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n157) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U155 ( 
        .A1(CurSAD[9]), .A2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n140), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n191) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U154 ( 
        .B1(extimating_unit_Results_calculator_SAD_min[8]), .B2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n152), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n191), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n195) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U153 ( 
        .A1(CurSAD[13]), .A2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n137), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n185) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U152 ( 
        .A1(CurSAD[15]), .A2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n136), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n187) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U151 ( 
        .B1(extimating_unit_Results_calculator_SAD_min[14]), .B2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n149), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n187), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n196) );
  OAI211_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U150 ( 
        .C1(extimating_unit_Results_calculator_SAD_min[12]), .C2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n150), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n185), .B(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n135), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n179) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U149 ( 
        .A1(CurSAD[11]), .A2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n139), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n193) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U148 ( 
        .B1(extimating_unit_Results_calculator_SAD_min[10]), .B2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n151), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n193), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n194) );
  NOR3_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U147 ( 
        .A1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n195), 
        .A2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n179), 
        .A3(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n194), 
        .ZN(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n159)
         );
  NAND3_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U146 ( 
        .A1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n193), 
        .A2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n151), 
        .A3(extimating_unit_Results_calculator_SAD_min[10]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n192) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U145 ( 
        .B1(CurSAD[11]), .B2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n139), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n192), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n188) );
  NAND3_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U144 ( 
        .A1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n191), 
        .A2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n152), 
        .A3(extimating_unit_Results_calculator_SAD_min[8]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n190) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U143 ( 
        .B1(CurSAD[9]), .B2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n140), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n190), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n189) );
  OAI22_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U142 ( 
        .A1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n138), 
        .A2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n188), 
        .B1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n188), 
        .B2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n189), 
        .ZN(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n180)
         );
  NAND3_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U141 ( 
        .A1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n187), 
        .A2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n149), 
        .A3(extimating_unit_Results_calculator_SAD_min[14]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n186) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U140 ( 
        .B1(CurSAD[15]), .B2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n136), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n186), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n182) );
  NAND3_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U139 ( 
        .A1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n185), 
        .A2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n150), 
        .A3(extimating_unit_Results_calculator_SAD_min[12]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n184) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U138 ( 
        .B1(CurSAD[13]), .B2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n137), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n184), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n183) );
  OAI22_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U137 ( 
        .A1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n135), 
        .A2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n182), 
        .B1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n182), 
        .B2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n183), 
        .ZN(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n181)
         );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U136 ( 
        .B1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n179), 
        .B2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n180), 
        .A(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n181), 
        .ZN(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n160)
         );
  NAND2_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U135 ( 
        .A1(CurSAD[3]), .A2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n146), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n178) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U134 ( 
        .B1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n155), 
        .B2(extimating_unit_Results_calculator_SAD_min[2]), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n178), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n172) );
  NAND3_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U133 ( 
        .A1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n178), 
        .A2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n155), 
        .A3(extimating_unit_Results_calculator_SAD_min[2]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n177) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U132 ( 
        .B1(CurSAD[3]), .B2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n146), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n177), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n174) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U131 ( 
        .A1(CurSAD[7]), .A2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n143), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n169) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U130 ( 
        .B1(extimating_unit_Results_calculator_SAD_min[6]), .B2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n153), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n169), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n170) );
  AOI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U129 ( 
        .B1(CurSAD[1]), .B2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n148), .A(
        CurSAD[0]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n176) );
  AOI22_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U128 ( 
        .A1(extimating_unit_Results_calculator_SAD_min[1]), .A2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n156), .B1(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n176), .B2(
        extimating_unit_Results_calculator_SAD_min[0]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n175) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U127 ( 
        .A1(CurSAD[5]), .A2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n144), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n167) );
  OAI221_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U126 ( 
        .B1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n147), 
        .B2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n174), 
        .C1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n154), 
        .C2(extimating_unit_Results_calculator_SAD_min[4]), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n167), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n173) );
  AOI211_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U125 ( 
        .C1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n172), 
        .C2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n145), 
        .A(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n170), 
        .B(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n173), 
        .ZN(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n171)
         );
  NAND3_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U124 ( 
        .A1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n169), 
        .A2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n153), 
        .A3(extimating_unit_Results_calculator_SAD_min[6]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n168) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U123 ( 
        .B1(CurSAD[7]), .B2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n143), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n168), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n164) );
  NAND3_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U122 ( 
        .A1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n167), 
        .A2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n154), 
        .A3(extimating_unit_Results_calculator_SAD_min[4]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n166) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U121 ( 
        .B1(CurSAD[5]), .B2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n144), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n166), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n165) );
  OAI22_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U120 ( 
        .A1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n142), 
        .A2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n164), 
        .B1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n164), 
        .B2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n165), 
        .ZN(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n163)
         );
  NAND2_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U119 ( 
        .A1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n141), 
        .A2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n163), 
        .ZN(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n161)
         );
  AOI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U118 ( 
        .B1(CurSAD[16]), .B2(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n134), .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n157), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n162) );
  OAI221_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U117 ( 
        .B1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n159), 
        .B2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n160), 
        .C1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n160), 
        .C2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n161), 
        .A(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n162), 
        .ZN(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n158)
         );
  OAI21_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U116 ( 
        .B1(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n132), 
        .B2(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n157), 
        .A(extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n158), 
        .ZN(extimating_unit_Results_calculator_ltmin) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U115 ( .A(
        extimating_unit_Results_calculator_SAD_min[1]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n148) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U114 ( .A(
        extimating_unit_Results_calculator_SAD_min[17]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n133) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U113 ( .A(
        extimating_unit_Results_calculator_SAD_min[13]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n137) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U112 ( .A(
        extimating_unit_Results_calculator_SAD_min[5]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n144) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U111 ( .A(
        extimating_unit_Results_calculator_SAD_min[15]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n136) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U110 ( .A(
        extimating_unit_Results_calculator_SAD_min[9]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n140) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U109 ( .A(
        extimating_unit_Results_calculator_SAD_min[11]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n139) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U108 ( .A(
        extimating_unit_Results_calculator_SAD_min[7]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n143) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U107 ( .A(
        extimating_unit_Results_calculator_SAD_min[3]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n146) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U106 ( .A(
        extimating_unit_Results_calculator_SAD_min[16]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n134) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U105 ( .A(
        CurSAD[1]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n156) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U104 ( .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n175), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n147) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U103 ( .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n196), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n135) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U102 ( .A(
        CurSAD[12]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n150) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U101 ( .A(
        CurSAD[4]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n154) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U100 ( .A(
        CurSAD[14]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n149) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U99 ( .A(
        CurSAD[8]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n152) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U98 ( .A(
        CurSAD[10]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n151) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U97 ( .A(
        CurSAD[6]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n153) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U96 ( .A(
        CurSAD[2]), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n155) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U95 ( .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n171), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n141) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U94 ( .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n197), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n132) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U93 ( .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n174), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n145) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U92 ( .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n194), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n138) );
  INV_X1 extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_U91 ( .A(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n170), .ZN(
        extimating_unit_Results_calculator_SAD_comparator_lt_gt_13_n142) );
  INV_X1 extimating_unit_Results_calculator_SAD_min_register_U41 ( .A(
        extimating_unit_Results_calculator_n202), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n58) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U40 ( .A1(
        CurSAD[17]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n54), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n18) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U39 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n36), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n57), .A(
        extimating_unit_Results_calculator_SAD_min_register_n18), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n55) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U38 ( .A1(
        CurSAD[16]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n54), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n17) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U37 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n35), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n57), .A(
        extimating_unit_Results_calculator_SAD_min_register_n17), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n53) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U36 ( .A1(
        CurSAD[15]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n54), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n16) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U35 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n34), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n57), .A(
        extimating_unit_Results_calculator_SAD_min_register_n16), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n52) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U34 ( .A1(
        CurSAD[14]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n54), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n15) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U33 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n33), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n57), .A(
        extimating_unit_Results_calculator_SAD_min_register_n15), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n51) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U32 ( .A1(
        CurSAD[13]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n54), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n14) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U31 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n32), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n57), .A(
        extimating_unit_Results_calculator_SAD_min_register_n14), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n50) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U30 ( .A1(
        CurSAD[12]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n54), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n13) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U29 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n31), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n57), .A(
        extimating_unit_Results_calculator_SAD_min_register_n13), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n49) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U28 ( .A1(
        CurSAD[11]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n54), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n12) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U27 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n30), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n56), .A(
        extimating_unit_Results_calculator_SAD_min_register_n12), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n48) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U26 ( .A1(
        CurSAD[10]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n54), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n11) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U25 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n29), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n56), .A(
        extimating_unit_Results_calculator_SAD_min_register_n11), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n47) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U24 ( .A1(
        CurSAD[9]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n54), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n10) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U23 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n28), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n56), .A(
        extimating_unit_Results_calculator_SAD_min_register_n10), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n46) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U22 ( .A1(
        CurSAD[8]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n54), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n9) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U21 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n27), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n56), .A(
        extimating_unit_Results_calculator_SAD_min_register_n9), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n45) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U20 ( .A1(
        CurSAD[7]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n54), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n8) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U19 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n26), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n56), .A(
        extimating_unit_Results_calculator_SAD_min_register_n8), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n44) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U18 ( .A1(
        CurSAD[6]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n54), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n7) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U17 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n25), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n56), .A(
        extimating_unit_Results_calculator_SAD_min_register_n7), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n43) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U16 ( .A1(
        CurSAD[5]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n56), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n6) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U15 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n24), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n57), .A(
        extimating_unit_Results_calculator_SAD_min_register_n6), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n42) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U14 ( .A1(
        CurSAD[4]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n56), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n5) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U13 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n23), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n56), .A(
        extimating_unit_Results_calculator_SAD_min_register_n5), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n41) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U12 ( .A1(
        CurSAD[3]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n56), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n4) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U11 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n22), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n57), .A(
        extimating_unit_Results_calculator_SAD_min_register_n4), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n40) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U10 ( .A1(
        CurSAD[2]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n56), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n3) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U9 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n21), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n57), .A(
        extimating_unit_Results_calculator_SAD_min_register_n3), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n39) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U8 ( .A1(
        CurSAD[1]), .A2(
        extimating_unit_Results_calculator_SAD_min_register_n56), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n2) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U7 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n20), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n57), .A(
        extimating_unit_Results_calculator_SAD_min_register_n2), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n38) );
  NAND2_X1 extimating_unit_Results_calculator_SAD_min_register_U6 ( .A1(
        extimating_unit_Results_calculator_SAD_min_register_n57), .A2(
        CurSAD[0]), .ZN(extimating_unit_Results_calculator_SAD_min_register_n1) );
  OAI21_X1 extimating_unit_Results_calculator_SAD_min_register_U5 ( .B1(
        extimating_unit_Results_calculator_SAD_min_register_n19), .B2(
        extimating_unit_Results_calculator_SAD_min_register_n57), .A(
        extimating_unit_Results_calculator_SAD_min_register_n1), .ZN(
        extimating_unit_Results_calculator_SAD_min_register_n37) );
  BUF_X1 extimating_unit_Results_calculator_SAD_min_register_U4 ( .A(
        extimating_unit_Results_calculator_Found_best), .Z(
        extimating_unit_Results_calculator_SAD_min_register_n57) );
  BUF_X1 extimating_unit_Results_calculator_SAD_min_register_U3 ( .A(
        extimating_unit_Results_calculator_Found_best), .Z(
        extimating_unit_Results_calculator_SAD_min_register_n56) );
  BUF_X1 extimating_unit_Results_calculator_SAD_min_register_U2 ( .A(
        extimating_unit_Results_calculator_Found_best), .Z(
        extimating_unit_Results_calculator_SAD_min_register_n54) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_6_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n43), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[6]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n25) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_7_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n44), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[7]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n26) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_8_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n45), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[8]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n27) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_9_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n46), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[9]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n28) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_10_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n47), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[10]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n29) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_11_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n48), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[11]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n30) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_12_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n49), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[12]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n31) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_13_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n50), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[13]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n32) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_14_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n51), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[14]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n33) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_15_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n52), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[15]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n34) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_16_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n53), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[16]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n35) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_17_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n55), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[17]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n36) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_4_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n41), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[4]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n23) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_1_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n38), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[1]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n20) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_2_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n39), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[2]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n21) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_3_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n40), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[3]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n22) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_5_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n42), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[5]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n24) );
  DFFS_X1 extimating_unit_Results_calculator_SAD_min_register_Q_int_reg_0_ ( 
        .D(extimating_unit_Results_calculator_SAD_min_register_n37), .CK(clk), 
        .SN(extimating_unit_Results_calculator_SAD_min_register_n58), .Q(
        extimating_unit_Results_calculator_SAD_min[0]), .QN(
        extimating_unit_Results_calculator_SAD_min_register_n19) );
  INV_X1 extimating_unit_Results_calculator_CurCand_counter_U2 ( .A(
        extimating_unit_Results_calculator_n203), .ZN(
        extimating_unit_Results_calculator_CurCand_counter_n1) );
  DFFR_X1 extimating_unit_Results_calculator_CurCand_counter_Q_int_reg ( .D(
        extimating_unit_Results_calculator_CurCand_counter_n2), .CK(clk), .RN(
        extimating_unit_Results_calculator_CurCand_counter_n1), .Q(
        extimating_unit_Results_calculator_CurCand) );
  XOR2_X1 extimating_unit_Results_calculator_CurCand_counter_U3 ( .A(
        extimating_unit_Results_calculator_CurCand), .B(eComp_EN), .Z(
        extimating_unit_Results_calculator_CurCand_counter_n2) );
  INV_X1 extimating_unit_Results_calculator_BestCand_register_U4 ( .A(
        extimating_unit_Results_calculator_n203), .ZN(
        extimating_unit_Results_calculator_BestCand_register_n3) );
  NAND2_X1 extimating_unit_Results_calculator_BestCand_register_U3 ( .A1(
        extimating_unit_Results_calculator_Found_best), .A2(
        extimating_unit_Results_calculator_CurCand), .ZN(
        extimating_unit_Results_calculator_BestCand_register_n1) );
  OAI21_X1 extimating_unit_Results_calculator_BestCand_register_U2 ( .B1(
        extimating_unit_Results_calculator_BestCand_register_n2), .B2(
        extimating_unit_Results_calculator_Found_best), .A(
        extimating_unit_Results_calculator_BestCand_register_n1), .ZN(
        extimating_unit_Results_calculator_BestCand_register_n4) );
  DFFR_X1 extimating_unit_Results_calculator_BestCand_register_Q_int_reg ( .D(
        extimating_unit_Results_calculator_BestCand_register_n4), .CK(clk), 
        .RN(extimating_unit_Results_calculator_BestCand_register_n3), .Q(
        BestCand), .QN(extimating_unit_Results_calculator_BestCand_register_n2) );
  XOR2_X1 extimating_unit_Results_calculator_Terminal_counter_U16 ( .A(
        extimating_unit_Results_calculator_Terminal_counter_add_23_carry[4]), 
        .B(extimating_unit_Results_calculator_Terminal_counter_count_4_), .Z(
        extimating_unit_Results_calculator_Terminal_counter_N6) );
  INV_X1 extimating_unit_Results_calculator_Terminal_counter_U15 ( .A(
        extimating_unit_Results_calculator_n203), .ZN(
        extimating_unit_Results_calculator_Terminal_counter_n7) );
  NOR3_X1 extimating_unit_Results_calculator_Terminal_counter_U14 ( .A1(
        extimating_unit_Results_calculator_Terminal_counter_n11), .A2(
        extimating_unit_Results_calculator_Terminal_counter_n8), .A3(
        extimating_unit_Results_calculator_Terminal_counter_count_0_), .ZN(
        extimating_unit_Results_calculator_Terminal_counter_n6) );
  AND3_X1 extimating_unit_Results_calculator_Terminal_counter_U13 ( .A1(
        extimating_unit_Results_calculator_Terminal_counter_n6), .A2(
        extimating_unit_Results_calculator_Terminal_counter_n10), .A3(
        extimating_unit_Results_calculator_Terminal_counter_n9), .ZN(
        CountTerm_OUT) );
  NAND2_X1 extimating_unit_Results_calculator_Terminal_counter_U12 ( .A1(
        extimating_unit_Results_calculator_Terminal_counter_N2), .A2(
        CountTerm_EN), .ZN(
        extimating_unit_Results_calculator_Terminal_counter_n5) );
  OAI21_X1 extimating_unit_Results_calculator_Terminal_counter_U11 ( .B1(
        extimating_unit_Results_calculator_Terminal_counter_N2), .B2(
        CountTerm_EN), .A(
        extimating_unit_Results_calculator_Terminal_counter_n5), .ZN(
        extimating_unit_Results_calculator_Terminal_counter_n18) );
  NAND2_X1 extimating_unit_Results_calculator_Terminal_counter_U10 ( .A1(
        extimating_unit_Results_calculator_Terminal_counter_N3), .A2(
        CountTerm_EN), .ZN(
        extimating_unit_Results_calculator_Terminal_counter_n4) );
  OAI21_X1 extimating_unit_Results_calculator_Terminal_counter_U9 ( .B1(
        extimating_unit_Results_calculator_Terminal_counter_n11), .B2(
        CountTerm_EN), .A(
        extimating_unit_Results_calculator_Terminal_counter_n4), .ZN(
        extimating_unit_Results_calculator_Terminal_counter_n16) );
  NAND2_X1 extimating_unit_Results_calculator_Terminal_counter_U8 ( .A1(
        extimating_unit_Results_calculator_Terminal_counter_N4), .A2(
        CountTerm_EN), .ZN(
        extimating_unit_Results_calculator_Terminal_counter_n3) );
  OAI21_X1 extimating_unit_Results_calculator_Terminal_counter_U7 ( .B1(
        extimating_unit_Results_calculator_Terminal_counter_n10), .B2(
        CountTerm_EN), .A(
        extimating_unit_Results_calculator_Terminal_counter_n3), .ZN(
        extimating_unit_Results_calculator_Terminal_counter_n15) );
  NAND2_X1 extimating_unit_Results_calculator_Terminal_counter_U6 ( .A1(
        extimating_unit_Results_calculator_Terminal_counter_N5), .A2(
        CountTerm_EN), .ZN(
        extimating_unit_Results_calculator_Terminal_counter_n2) );
  OAI21_X1 extimating_unit_Results_calculator_Terminal_counter_U5 ( .B1(
        extimating_unit_Results_calculator_Terminal_counter_n9), .B2(
        CountTerm_EN), .A(
        extimating_unit_Results_calculator_Terminal_counter_n2), .ZN(
        extimating_unit_Results_calculator_Terminal_counter_n14) );
  NAND2_X1 extimating_unit_Results_calculator_Terminal_counter_U4 ( .A1(
        extimating_unit_Results_calculator_Terminal_counter_N6), .A2(
        CountTerm_EN), .ZN(
        extimating_unit_Results_calculator_Terminal_counter_n1) );
  OAI21_X1 extimating_unit_Results_calculator_Terminal_counter_U3 ( .B1(
        extimating_unit_Results_calculator_Terminal_counter_n8), .B2(
        CountTerm_EN), .A(
        extimating_unit_Results_calculator_Terminal_counter_n1), .ZN(
        extimating_unit_Results_calculator_Terminal_counter_n13) );
  DFFR_X1 extimating_unit_Results_calculator_Terminal_counter_count_reg_4_ ( 
        .D(extimating_unit_Results_calculator_Terminal_counter_n13), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Terminal_counter_n7), .Q(
        extimating_unit_Results_calculator_Terminal_counter_count_4_), .QN(
        extimating_unit_Results_calculator_Terminal_counter_n8) );
  DFFR_X1 extimating_unit_Results_calculator_Terminal_counter_count_reg_0_ ( 
        .D(extimating_unit_Results_calculator_Terminal_counter_n18), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Terminal_counter_n7), .Q(
        extimating_unit_Results_calculator_Terminal_counter_count_0_), .QN(
        extimating_unit_Results_calculator_Terminal_counter_N2) );
  DFFR_X1 extimating_unit_Results_calculator_Terminal_counter_count_reg_1_ ( 
        .D(extimating_unit_Results_calculator_Terminal_counter_n16), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Terminal_counter_n7), .Q(
        extimating_unit_Results_calculator_Terminal_counter_count_1_), .QN(
        extimating_unit_Results_calculator_Terminal_counter_n11) );
  DFFR_X1 extimating_unit_Results_calculator_Terminal_counter_count_reg_2_ ( 
        .D(extimating_unit_Results_calculator_Terminal_counter_n15), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Terminal_counter_n7), .Q(
        extimating_unit_Results_calculator_Terminal_counter_count_2_), .QN(
        extimating_unit_Results_calculator_Terminal_counter_n10) );
  DFFR_X1 extimating_unit_Results_calculator_Terminal_counter_count_reg_3_ ( 
        .D(extimating_unit_Results_calculator_Terminal_counter_n14), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Terminal_counter_n7), .Q(
        extimating_unit_Results_calculator_Terminal_counter_count_3_), .QN(
        extimating_unit_Results_calculator_Terminal_counter_n9) );
  HA_X1 extimating_unit_Results_calculator_Terminal_counter_add_23_U1_1_3 ( 
        .A(extimating_unit_Results_calculator_Terminal_counter_count_3_), .B(
        extimating_unit_Results_calculator_Terminal_counter_add_23_carry[3]), 
        .CO(
        extimating_unit_Results_calculator_Terminal_counter_add_23_carry[4]), 
        .S(extimating_unit_Results_calculator_Terminal_counter_N5) );
  HA_X1 extimating_unit_Results_calculator_Terminal_counter_add_23_U1_1_2 ( 
        .A(extimating_unit_Results_calculator_Terminal_counter_count_2_), .B(
        extimating_unit_Results_calculator_Terminal_counter_add_23_carry[2]), 
        .CO(
        extimating_unit_Results_calculator_Terminal_counter_add_23_carry[3]), 
        .S(extimating_unit_Results_calculator_Terminal_counter_N4) );
  HA_X1 extimating_unit_Results_calculator_Terminal_counter_add_23_U1_1_1 ( 
        .A(extimating_unit_Results_calculator_Terminal_counter_count_1_), .B(
        extimating_unit_Results_calculator_Terminal_counter_count_0_), .CO(
        extimating_unit_Results_calculator_Terminal_counter_add_23_carry[2]), 
        .S(extimating_unit_Results_calculator_Terminal_counter_N3) );
  INV_X1 extimating_unit_Results_calculator_Candidate_counter_U2 ( .A(
        extimating_unit_RST2_int), .ZN(
        extimating_unit_Results_calculator_Candidate_counter_n1) );
  XOR2_X1 extimating_unit_Results_calculator_Candidate_counter_U3 ( .A(
        last_cand), .B(ADD3_MVin_LE_nSET), .Z(
        extimating_unit_Results_calculator_Candidate_counter_n3) );
  DFFR_X1 extimating_unit_Results_calculator_Candidate_counter_Q_int_reg ( .D(
        extimating_unit_Results_calculator_Candidate_counter_n3), .CK(clk), 
        .RN(extimating_unit_Results_calculator_Candidate_counter_n1), .Q(
        last_cand) );
  XOR2_X1 extimating_unit_Results_calculator_add_85_U17 ( .A(
        extimating_unit_Results_calculator_SAD_tmp[0]), .B(
        extimating_unit_Results_calculator_CurRowSAD[0]), .Z(
        extimating_unit_Results_calculator_CurSAD_tmp_0_) );
  NAND2_X1 extimating_unit_Results_calculator_add_85_U16 ( .A1(
        extimating_unit_Results_calculator_SAD_tmp[16]), .A2(
        extimating_unit_Results_calculator_add_85_n6), .ZN(
        extimating_unit_Results_calculator_add_85_n17) );
  XNOR2_X1 extimating_unit_Results_calculator_add_85_U15 ( .A(
        extimating_unit_Results_calculator_SAD_tmp[17]), .B(
        extimating_unit_Results_calculator_add_85_n17), .ZN(
        extimating_unit_Results_calculator_CurSAD_tmp_17_) );
  XOR2_X1 extimating_unit_Results_calculator_add_85_U14 ( .A(
        extimating_unit_Results_calculator_SAD_tmp[16]), .B(
        extimating_unit_Results_calculator_add_85_n6), .Z(
        extimating_unit_Results_calculator_CurSAD_tmp_16_) );
  XOR2_X1 extimating_unit_Results_calculator_add_85_U13 ( .A(
        extimating_unit_Results_calculator_SAD_tmp[15]), .B(
        extimating_unit_Results_calculator_add_85_n5), .Z(
        extimating_unit_Results_calculator_CurSAD_tmp_15_) );
  XOR2_X1 extimating_unit_Results_calculator_add_85_U12 ( .A(
        extimating_unit_Results_calculator_SAD_tmp[14]), .B(
        extimating_unit_Results_calculator_add_85_n4), .Z(
        extimating_unit_Results_calculator_CurSAD_tmp_14_) );
  XOR2_X1 extimating_unit_Results_calculator_add_85_U11 ( .A(
        extimating_unit_Results_calculator_SAD_tmp[13]), .B(
        extimating_unit_Results_calculator_add_85_n3), .Z(
        extimating_unit_Results_calculator_CurSAD_tmp_13_) );
  XOR2_X1 extimating_unit_Results_calculator_add_85_U10 ( .A(
        extimating_unit_Results_calculator_SAD_tmp[12]), .B(
        extimating_unit_Results_calculator_add_85_n2), .Z(
        extimating_unit_Results_calculator_CurSAD_tmp_12_) );
  XOR2_X1 extimating_unit_Results_calculator_add_85_U9 ( .A(
        extimating_unit_Results_calculator_SAD_tmp[11]), .B(
        extimating_unit_Results_calculator_add_85_n1), .Z(
        extimating_unit_Results_calculator_CurSAD_tmp_11_) );
  XOR2_X1 extimating_unit_Results_calculator_add_85_U8 ( .A(
        extimating_unit_Results_calculator_SAD_tmp[10]), .B(
        extimating_unit_Results_calculator_add_85_carry_10_), .Z(
        extimating_unit_Results_calculator_CurSAD_tmp_10_) );
  AND2_X1 extimating_unit_Results_calculator_add_85_U7 ( .A1(
        extimating_unit_Results_calculator_SAD_tmp[0]), .A2(
        extimating_unit_Results_calculator_CurRowSAD[0]), .ZN(
        extimating_unit_Results_calculator_add_85_n7) );
  AND2_X1 extimating_unit_Results_calculator_add_85_U6 ( .A1(
        extimating_unit_Results_calculator_SAD_tmp[15]), .A2(
        extimating_unit_Results_calculator_add_85_n5), .ZN(
        extimating_unit_Results_calculator_add_85_n6) );
  AND2_X1 extimating_unit_Results_calculator_add_85_U5 ( .A1(
        extimating_unit_Results_calculator_SAD_tmp[14]), .A2(
        extimating_unit_Results_calculator_add_85_n4), .ZN(
        extimating_unit_Results_calculator_add_85_n5) );
  AND2_X1 extimating_unit_Results_calculator_add_85_U4 ( .A1(
        extimating_unit_Results_calculator_SAD_tmp[13]), .A2(
        extimating_unit_Results_calculator_add_85_n3), .ZN(
        extimating_unit_Results_calculator_add_85_n4) );
  AND2_X1 extimating_unit_Results_calculator_add_85_U3 ( .A1(
        extimating_unit_Results_calculator_SAD_tmp[12]), .A2(
        extimating_unit_Results_calculator_add_85_n2), .ZN(
        extimating_unit_Results_calculator_add_85_n3) );
  AND2_X1 extimating_unit_Results_calculator_add_85_U2 ( .A1(
        extimating_unit_Results_calculator_SAD_tmp[11]), .A2(
        extimating_unit_Results_calculator_add_85_n1), .ZN(
        extimating_unit_Results_calculator_add_85_n2) );
  AND2_X1 extimating_unit_Results_calculator_add_85_U1 ( .A1(
        extimating_unit_Results_calculator_SAD_tmp[10]), .A2(
        extimating_unit_Results_calculator_add_85_carry_10_), .ZN(
        extimating_unit_Results_calculator_add_85_n1) );
  FA_X1 extimating_unit_Results_calculator_add_85_U1_1 ( .A(
        extimating_unit_Results_calculator_CurRowSAD[1]), .B(
        extimating_unit_Results_calculator_SAD_tmp[1]), .CI(
        extimating_unit_Results_calculator_add_85_n7), .CO(
        extimating_unit_Results_calculator_add_85_carry_2_), .S(
        extimating_unit_Results_calculator_CurSAD_tmp_1_) );
  FA_X1 extimating_unit_Results_calculator_add_85_U1_2 ( .A(
        extimating_unit_Results_calculator_CurRowSAD[2]), .B(
        extimating_unit_Results_calculator_SAD_tmp[2]), .CI(
        extimating_unit_Results_calculator_add_85_carry_2_), .CO(
        extimating_unit_Results_calculator_add_85_carry_3_), .S(
        extimating_unit_Results_calculator_CurSAD_tmp_2_) );
  FA_X1 extimating_unit_Results_calculator_add_85_U1_3 ( .A(
        extimating_unit_Results_calculator_CurRowSAD[3]), .B(
        extimating_unit_Results_calculator_SAD_tmp[3]), .CI(
        extimating_unit_Results_calculator_add_85_carry_3_), .CO(
        extimating_unit_Results_calculator_add_85_carry_4_), .S(
        extimating_unit_Results_calculator_CurSAD_tmp_3_) );
  FA_X1 extimating_unit_Results_calculator_add_85_U1_4 ( .A(
        extimating_unit_Results_calculator_CurRowSAD[4]), .B(
        extimating_unit_Results_calculator_SAD_tmp[4]), .CI(
        extimating_unit_Results_calculator_add_85_carry_4_), .CO(
        extimating_unit_Results_calculator_add_85_carry_5_), .S(
        extimating_unit_Results_calculator_CurSAD_tmp_4_) );
  FA_X1 extimating_unit_Results_calculator_add_85_U1_5 ( .A(
        extimating_unit_Results_calculator_CurRowSAD[5]), .B(
        extimating_unit_Results_calculator_SAD_tmp[5]), .CI(
        extimating_unit_Results_calculator_add_85_carry_5_), .CO(
        extimating_unit_Results_calculator_add_85_carry_6_), .S(
        extimating_unit_Results_calculator_CurSAD_tmp_5_) );
  FA_X1 extimating_unit_Results_calculator_add_85_U1_6 ( .A(
        extimating_unit_Results_calculator_CurRowSAD[6]), .B(
        extimating_unit_Results_calculator_SAD_tmp[6]), .CI(
        extimating_unit_Results_calculator_add_85_carry_6_), .CO(
        extimating_unit_Results_calculator_add_85_carry_7_), .S(
        extimating_unit_Results_calculator_CurSAD_tmp_6_) );
  FA_X1 extimating_unit_Results_calculator_add_85_U1_7 ( .A(
        extimating_unit_Results_calculator_CurRowSAD[7]), .B(
        extimating_unit_Results_calculator_SAD_tmp[7]), .CI(
        extimating_unit_Results_calculator_add_85_carry_7_), .CO(
        extimating_unit_Results_calculator_add_85_carry_8_), .S(
        extimating_unit_Results_calculator_CurSAD_tmp_7_) );
  FA_X1 extimating_unit_Results_calculator_add_85_U1_8 ( .A(
        extimating_unit_Results_calculator_CurRowSAD[8]), .B(
        extimating_unit_Results_calculator_SAD_tmp[8]), .CI(
        extimating_unit_Results_calculator_add_85_carry_8_), .CO(
        extimating_unit_Results_calculator_add_85_carry_9_), .S(
        extimating_unit_Results_calculator_CurSAD_tmp_8_) );
  FA_X1 extimating_unit_Results_calculator_add_85_U1_9 ( .A(
        extimating_unit_Results_calculator_CurRowSAD[9]), .B(
        extimating_unit_Results_calculator_SAD_tmp[9]), .CI(
        extimating_unit_Results_calculator_add_85_carry_9_), .CO(
        extimating_unit_Results_calculator_add_85_carry_10_), .S(
        extimating_unit_Results_calculator_CurSAD_tmp_9_) );
endmodule

